-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OdJ6mIUqPJDYwSQ0lE3vpHKHYv5Hyzmz0d1I89QXQXJU8L4kgnw8I1ibTIoWfyrc7WA6Q3b5TgGg
ntSd9gmwxM8x2GB4FvH0M9e6m4rfOYkuk11Qa4Ozfw/XvEAt3zDQT7wrPj16km/jXl7og09d2b6c
501YsRmx3fw8sY01QijDj4T7ur5dy6W5Mpk5iyWXH6Uf02M2WkdamQoI9VzNhAH12XJ/twxNDRw7
Oqq/pVb9I4CuCEEy9BdjpuPbkvAJ5DHBTBEt6PvWcBGCxwHQMy73/0pSSBx5Dv/cYUH/18P+Zo5h
7N7tFc/szkzDe5YluFSJLoBvIBULIFlRuPJP9Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28512)
`protect data_block
uGdNG4bHcQP2VPQL2xZuVmIPSqhydwsknD6k6y6jReFwxwu1YLz1CKbkfpY7eXgPkEagNFvhygJj
azsRyITgc09emM0MrCFXuj5WSc9QHToNd+ucNcYGaG944q6L0FIoWo4R/7vjCfH49MQDh+O+ULJ7
263tkY9kL/Cm75k52NmvqSFAIPNRiStUt84wiy+gA82+WkxQ3m6XikJ3ql/GDdVMHdzw0mqUUIPD
B/boVTQSQc6ucKiktjhouggB3xG2w9pPINOC97V7A7TZYKtMPmrsXKq3NMFoej4Jk1sk5pvp6Xy8
QB14XF/ucGvBvv/jIa9FGdla0uIXDGuPOlEVawsgqfgr0K7Qb4X8TiEV0tkBcTpjSMBD1SEt6NuO
WvU6k8qljUMPwyH3AttyxZ7K8KBPYWT+KcY00k8GZYPxSkV/+m6ZQuTV7/Dzza/pgZKipLTPkDfa
lWrJkks5kETDyF0QM2a7RkemUKwqdbtGxY0js+1GyALi9r0xD20WIkrL+gNFE/mBaK9RYxkKejPX
u1LGVj451CYNmi4ELstljczgsjE2xR2KWbcQB3Lz9mxce86eiODSuNlcfSmM6PhPcv8C/iuEigdN
pUH2iPmaQ/p+Rm35vXiM6UUmTb0vMVBE4BKgWQfdgQdqBLZRmGCKhqLfpdNllic7ZCQLG1L7iUan
lnREHwVpuJzm7M22u/Xw/Yi8E710/xQg4ZHqTD93ri0S3gUaYNy9qUg5LMy9xwu/+Tdgiz5ZbCYz
+gWBqxqomQ9mAAQwP3XTJNoyqbnBz/z3JF+SjxrTVYi1JSLuWHvM0oTnzuazgm7sOiJARe+fYR8c
UpX8rRE46eXCtyPaa6Y5DwkVrUjljBwS4cYSfqQwcDc/+Nh/dw9zkxa32IOqJizs3vVA10khW6wA
7imLh5K7pDhINRTGKy84Mb3UTNehb2FBghnxsIrp8BZ0Gi20lDe2vESwy1z3v0LlCZJumjTfkOOF
PXZTBz57XaiGtUKNrxKExt1EhPC25gfLVRrfN5gHpW+ti0HgdzqxrQDdH4gkxvsh6srGF5uH1HF4
MKOJ6PqclI4+HhtmsbNWFvVyfPIDz6NTEUWtLjokWGSTkYDpHip8CKV2iFYSZcDABvrbN7vyjmva
WlOV9DaHx/XwiOlHTHBTMdDVbaubsQ2YFOzaZ5tLJwBAMnMGXbzd8i/CLLWFguS+Afxbvs8xCj5f
x0GxmUvMsOsk1IQCHrRYXIOl+7XIhzKxHM/eRePzu1MHWsP+9vcIIshb1DgUbV0c+cRnzIIMz2MA
KJKpYfnesVtv0ZRBjbiqd9NGT4l019YiyD9C/nMcBj+WWCfiJEnjJbGnBvXaQsKKRkhkH2ShFOaI
SECjTZxGne3bUB/6NLzn6Whq61ZW635YysjnS2pwqcING8yhHnMVuocFV4i8uIHBPpqXE/59oEKm
DxVaaWYxNWMIkZTzPvjS1bSoelOOq0IyKguM8tl+aIlw55brpvs/1sRcI3L03Op32FG646iicUHz
QzTCPpZq5wXjpGiCyM4COIyt8b8N3MQ0NayeDR5845R/mD/Dl6EYutf5CuiW3lAnyTL9xlW2Hx2A
gcmdewER/bHHa4F0Eme11SqL9DTvoCvJboMA9GaE1OP+gqqSJWLTNO4KqQZCvy6qtjDcpZp2Mniy
fdp7VavitDzf8RcOGyW5URzxC/6X9A6aqyrfjrDn7DiaJCkoFz7v6gQ45e5sPup9B3ewq8iXGCXy
11y/BWvJg6iG3MU5LV9uXb2kIIrcaodmyo+gtDd+SwC9ajPn+EiTSpDAWLA6iFSoqto1KKlydCml
Qd9t2qgA0tkXLbzvtBaPxR+94PHkgWTd4BZgq65SM9u1gBw0F/TgQW4F4fZJqle/RipxYwPszbEh
xwZ9asxZx8gINH22B1oYRC371fjNeUZh1BGxr54nXDc5QQ7e1ZkLDwhA/eU9D1Ab6kbxLR2EBcRD
APghvxA9L2o5Kx8HES+ZRaFoEwTkRjYj9dglK+/IqCJujassGIC2JpHRQlPDtNCqrcid4hLMmdct
XmFwen1HQq0XyrVtiNMVABVmka2bnRySYQXHo5vin7DnBOyms74VUArVa15C4NNxu/ulVhq7MUrZ
pF4joLZskHwOmTj0y9DRGxxPM3oVnNTd5ZkQlrlGDB6XYtdtEK7yKGA6WJGfhdtJjpU8QHpZiJgX
GNnVq5q5t4eB0g9ccpjg8rfLoiO15aV+Tkp/GoukVYj7h0tn/gsml0sFU3+znuXJN/D5eiajs1be
djM6A2k4p6jFrVUVCdhxdIE8q3uO3obdvbdEo6OiB0zHmM3cZf41zR++CwdJ6JucdmgXAGQmyp8u
NNHAtbsOFt6GnUpTE+HEWoZJc88KlsulWw3wABLmQNphf4ER2Lt0KNJiCFuRB37Zapj46w4oRNe3
Z/Fd5/e5Z9v5rFgA+661au5jli3k8gjk07XdIUadK5ho9xZsQMUdR6nENtw1kHlKPrM5RfwW9h1+
uxWe0taUxXEdJSPeDUzMeSOHpIFpk40PIbYUUwoP+Li6sKf55p3XMdeCddXn59iJz1NkJeSPJN/+
Xci8SE80iCBC6tSij+5BpsBs7C7LOzPVdfvE+JP2lQgB7L9kywAlmZi3XtqAKS0JG4aQA9mEkrYw
P4HtDWNfAcMbWd57I4HjeizB9nkPsMtzzKVtiL7Xse2vgmH+cdEuj12of4D9oTT5HoeQ/eSY48Hm
iljjtZq95HxlKTXQkc/W/Pp9OuGKhS9UOsyw5q8GzYL3t1oB65IH/4Pg7vNFUOt6PVAsfiu9jwEx
J+adlbgJ5E0Dw5BOndgVHapnzAyfe4Cdh7NWqyLypWbk97LGdw7CfHgNgyp5keea38Uy3Us45MwY
Jn3nGv2m7VJkEZtDmD4BRQKwlRS9jNYJatYltXBnVSCvQbM+fCst/wRMuoDX447RqXXHz/3IHM5b
qzYZgAduk8NgSK4zI48oiyi/H1OHpLB8OTckw6VYwjXddoFMZZZZR0WqpLmeQWE/yioJdw0SRD0o
2CXErVnO/rRqKOMDSoLQ8+cC3fZwPxNRH6YtNh9yEgPp2BghaIwSTtZT8eCcnubeY+i4Me1Kj1dE
NLTkl/xQsd7h25ZpDvPNbjBgEFewBvBdup1LxiWWB5ZDmcN7IfuJTaT7czx7q4lB/EZq+R2NkeJh
oDYEGS0vlRdukZAWYY52JjGhqLvQzIXKBc0T5/+5gx9m8s0D9LQtq8TodoQX3IORKO5AZ9YYO590
431haAmNweD4zCPKafVgSi5kDZPuxUZX+lv5sdkjee2oG08AvpVeY9ZbriQH4IMAvH6sJ/Hl/Vxq
kpWVQdO3g6cSckswHui6K7qsSDYSeNH+3gsZeVPROpqGp9wEkV/tCfjWUWMJK8Q2F07iG0ZCg0k2
74W14Rwf9K8lDJMHauchceaH8n8H16+Q6tqQbf/wdx6wpYNYYWqw6kCTYQxzz3hh1a4SUKG8K2wj
Xl/plMaaHMMd83WxxTXehrR/KvYUSQqoy7Z6sxkrIjO7cq9BpUCwkjU8dTjZcQIxiw9NCp25+bWq
lAhZS2Lqb0mRS236sPUUqJ3E7xfc0yCOkT0n3Mwc/VhoiEy7C6FhkzWezNyb9dYyqXLgXm+6Q3PD
xct2rtQlpIzPa2LuasLCWxA3lgz2BxAbxvY/dbbDEg1S5nHQkqLoSYIXSlL2Q/05mU12Ro0HbtwX
mDJmd6RPz5bng00exKwtQ3Y8MiSMURE32c1iMoMvR4leevWE+kiuQw6+ROwMXtTZEU1cEzQK9p+A
8ec+OO84KcwXR84WShNP4DkSJJY2HDRPkMoLyaKhL0PrHl1qATYXe/P6GZd0u2DbS9ABeeSofeb4
AmtKK3dd2dc47ll4gaWhC0gu6UEaaaWtKqc/aX8LIqEIvx5Xucm/BhIPtAr0c/z+ATuP/nDXwofB
yj+ilgVN5htShMCVAvs2KgsxBVgslL/tJNgwnRUC6TUhDdDuYpEVGKFhy7C1nfVcOWuDHT16LHh0
xx2U2nr6C7zVQNwPZUNbsjWTynRShKcSYeTMD4uIQZ/8FGuoh32r1HmQxPP+Xp+q28bB2hmKg+HV
Nyj+GuakHgHM+y8uKI9PjYqVGjpXFMTWtZ4W6hg2cBi21b4tdBO0XbWp9Ljawq8+Ojot36FERqU2
aCzIN+zfp5AEpWnEi7HXsyA8/H5PE7FtZDJjrgs56uXxvFq6RC+J2RkYInzuhduuPPRQM3CtMnDX
EMtDd7R0edyH31iXFI9KGP770E+j0men4JUpEU417w6pKxhxtKnrw6fU7JEnKGq3qgAAB3JjVDMG
am7Z0QH2xtKWFYkJEqztMmsWOqVoUzritUj2/CwxqqbLBXChb0kBBBO5GCII7qsGX7c2IhUqcwqW
UIXYn1pHTHbNrCrIU6CKsaTQYPH/x/wRIG0ASLh3PcMtc6XtZnijCXgUmerVx0t0x1tF2iMwywI5
+zR0OoLeQ1b4fxlIJdhMqG7JrWQ3bWLlcFAzDlNHTf+GCqVp9Z4+jDvTRmaYADzVDcvJVp5TqYco
5tT6DsUO/WSm9ZjIlfQLHxB1QPEKvZgXX3XKwxx0khEoXCfGMws6HCed1l8O1YAuMOmb7A4JMKDl
vI/aEcs6b32vuHXPrp1+3KUE44jZPyx7nttaSGklsQJ6rbG5PlbqvimwKFL9N9QZ3bbR/T6MWAQX
/WslSdgf4yStVlusLeypIKIKhmwCOZeuvTSzZE+hbDZykII3olbfZwYlt0rgGPyDyXhVUxtQvZUC
yZF3/M3qiNNyTJG7tUwCJQkLEOrKGFR3TMV3Quio4aabyNCBkLb4vvQMNMDxl9ULhtdBmrOCNzjJ
ds7lhM0xJKxTv2b+M1osZTUxz3T/TLu03VaxFKKjjWgBYwv3KoxvzQ+ajBvByRkt9IuDTjkIMO0A
tBvWigFeqeR4M2G3OCXaxjV+0NbEpsNA7FOVXyKvYYfd9j+sDJIE8FLvtFR/7388I7bwgoQ9emXZ
oPjInj9EprACunBv25D5ecVzKpYbPa8CIXaiGLBUfzC85xDw0UWwx4ikfbTNeVfGpCjqp0C++j59
6YHwMXvZmpaTuHZXrtS1Zs+ld8RW8ls9uCEv+uuLD9Rai8vyIqWJL9WgsuBYgdR8mYplYfoa/PMc
AljM7g0qyqd/QARhmASRRAPJe6vkJ8/2YIYaisPQQgmzYq6HH1TFFrWHyGMiVe3SxvPLsuwHy9i+
6iShBWmU4YM87EvA5FeM4nMHrD9veObwF03UMvigAvJ5pF9fGwF3qebu/AOPEOcuO7BP7hjY8Gfk
zEPpRuVvjzDgliMro8iTWWYcmN2OgSd7/1PMwULdic+zO+oAQUrHS8jVWG27wh82CVtvqPpSw67H
OHDTxGwJyCChtExyO8Ln9UTqyf/axwxnAADe6VGaq9iLZAm3Gn3Mms6Iok3HVRZhc8XGpqq8bbrM
UmQW8Y7MAt75R1UaJxM5j1DaiPIwbMFyF6pSEzLIs6bjU7Cb1pWj/w7egvBJXtggRjzhrimUluuq
aUh75BrmURsknN7vFLGds5Jh/JL9T1KiPiWFRuglUZfFDMbgz0OiUyxRW6Gk9nu1KqexDT3im5Kj
Yc5uLylBP/oms5sluxvIrb5ptBJ3jH4+eDhw/nYgb0AjqaXyOQz8029QMCrKKD5luc+p9aFhXSmB
20A8/JzakNRm40XHrJK1MZpCjaC/GqDl+G4bYQwp+QahSdErv+rnvCL3aHQHfsfl47nkQIdPZqVJ
lUxCwAqXvLk9Ygc5kw497d+Duk/9M1qLjNy9FwuzRQIwP85SEWqvnI4SEVYtoDvKJWO7GXfUwmNf
v6aaqVKuL3HBGNVJkQ5QPWCmglz5RHUWBw/wqQKTyyJV6p3ONRmOYX00Y5e3+PheZvjxSHe6Pfce
3NES2AA43zJGDXFox+WpMLp2yqTDhLXINKz4a9LKGOMjrIkCoJcLu0M7F7cFd1gKvWmzy1xT+xYp
RoZOldgTxuGuAHhG9RQ3KwODxMH7s1wjqwrlHTLO9J5YSwiqWobY3xCEy4gZ1hCbdGe26V+iPdlk
kBpShLSMuH6MU+9W7yk6t2Stb6P6LL97SOCBXW9mVDF1iLPeYrIcza55fcuXVN7ZT5epJRLDoyQa
aOPKisbPWOrguhSjW3ej8G8wc8YV4HMiuDFmzA2YV/bGIrGl5PFRlHyI81RzIPRX1WCuQYFiZW72
rNPDHj6eU+sLqs5lxSkT2Jee8gPWiZxfxjKxB85py7hOOY7ac8oaCUaYpDrNkqKAhi7V3CDhjrGe
+53QCsl8Y7KFk7QX/RQw867qNeWfDYrHan7qaRQ6O1fme30UyUI+K4x8Jv5ZlAzyVjZME5eODTxq
ijl8Cuws0m1krU+CtP6KZ0w8XSJQdPXA85MkcMMvDqnsb1VSirk7Xkemqd6XF892CSzMXpRZnrdP
XnsjVha+TbZN2SDKzskNKtZSc9Cy94Gtjgsb1I16RCiLqFbNW/UzEPv0CxsQu6jS+d71tt3RFlhs
FouY9LSIsMTBP+ce35BZXDh4ppcrzKPdF/yTAoFuzj0km4JKzmFd/DcIPPFsW6ie8pHxksmupoh1
D9bCc8Ty0kECfjF7bsYRrGXS1RKl77S4/HANr5/UJAg5GBZX35BkPH97bItNuCAzxKK8GTkxrFsf
6UG9OGhYwSP4+rhSZWJhN4qeMSJJS7irxJG8fOI9qn08DDsT2H4vBAia0mcZ6rEIJRK9w/AycefL
A/8fdHRofIC1DOZaTMpXY6XELhOcFjqgIawClo4+y0QgGgJEuTSxknj2wIE92IAlaGYCBCufTC5U
ldQ7Iy0dzD4RN+pw+pN7P6/x3cqYzG3V+P96c4RLKG988az4/x66hsDE9SjFxKauoIZu94RTUmho
q5MDy5lfhZd5V70B69UVDQzN6285rzb/hQ1l8a34u+aE0OmBg5kPGtcxMZgTn83ATMYsylyMl53G
wxUKta+VV5qtiyj35f3/UBHnGKrHhIS/B/Ctwz8SmfK9dZo1F9WGeaJ02u19hMKeQ/+jvu74xW8L
cp+9lrHTHmmTWBsjWuFMlQ3UG2ag2VDT+SZYQe9u2GeQRn4mpcKRUYCF2maGYNv9v6ZKjou4hXM3
IokJZMfKXcxJbElxBFHRT/nz+RExJyCDj9gH8yC9iQ5uo22fHIjVw+jrLuBV/4YiV8W44ACoQq3r
9UKvUYtX0g/4XgOaHmQz0CCX1LwFoieyVu3jZm3AgVcvGYVdbRElTbblexyT8gcBb24RNNBZZo8x
QGAnlRDDERoMCbvFj2VJm/rU8f9o9rW21B8zGUl46sEjqrYr2bd4p+C0URt6bU7UCdHEuqNdD3ow
2e5+PCgZdd0WhSB6luUUKQAjXFyCc3ATB/OLD+L8QfgiBwYgnkRbPLTPM/xie/e1l5lZT6d2xaF+
0BAqkGKNuNW+cfmdtnf7p4kKOavJe6+pgmS98RzpCeITORg/xQvFX2/Lor5Jf89wXSIm/Gu7vrEU
bS/bGhnpgPKqK/W7AosoSIDW5onauc+P2aya/wUNiLPh7U6RV4QEipiCYgZphPRVDc/YTAewc9yx
WG/1F7UWnp93dE1YXSko5oiE9fBe/quoJM57yahnleif2WVjX6orjjDC/P/YwQpkeg1sKaZl/cKm
75PUD2Kis/lfOsdjs8M7KJuR7f8GWVI7ye8ZFO61/uDUN5LsOWr4bgvJf55hjtB3gVqu5Do5FfCm
eA8up0Ivvo3vdBRS6G7durES4N9EKGyEjHjc6jGMEUHGSgp6McTMabvOq1NmIPnzYzYn4z27py17
ZNH/eg9r7fmKex38NkssAIHnexQ8jNbvsouOcasgdPEQOrMNaFC2OfbO024jlCX8pFiu47q5vUrE
sJHwYdRmhS4caGC7X2u3igdINdVADdsz4/89cU/pYv58cOgIFMBe0B1bCLcJfr4F0JFh9kpN7PGe
0hXWFPVjIVKghFsyhMs5plcF6Bxk73Txt/KfsGuLeeztxdhAZnZzmdx4ToImn9Li0n1kCq4J8z68
enBu+ENJN6jhi+fn0/WR8byTOOEgPNSbA1JjG8x7jMPy2doX20sW8atvL80UsnYMr+wvK3Nw5gxx
G1yMvQxpJhjxWl4+ItuzRtD++OEKz9a6Cw0F9dhHI+i3jJsKZ6W42oOapv8lzxoC40gQydOwpZup
bYO2XQ1ltOPxbSG5dNB34cx9UJUvVBahMtnNiYicgldT5UuiLcjXnBqzcU7SDhwChgyJklTih2t1
e/8ntGlwgFML/x+T1jrlVKbip+geFuuc8mafIGZK1A+5X5M4y3lu8YKF70hV+pXedRtBd0oLBTSZ
/jSecMJqp+PfIfDyK+g8GnmwSpkWKIoJeMu5mpvCwR7trC9+om9WPZYMVl66VP0fpmoUhdyLOPIi
5Z9AAtgh+NqYR3rrCW+4kXBf0ltxmnV3ATxW7WHcnw9MLyzOdHcA1yx/f0gxKlTAzpF1+vYCaKSk
P3CbkIRvB7x8UZo4uS/Nk2gryO8R1xYnd2fMyXX6gu5Zndx3XcdudBepGVhUip0NOGrAFRoKDwBj
l9lzfQtzjE2ompTlUga9ONO9DS0PRUfS6DzUEWI9ovqYTkq06VddM+Kd4ZSpypI21ck7aRdH8bwp
z44MK1RE+mXsejPmRSQgkeanJkqup2cC/3ZsuyMJT63jtkpCNodAJmRAivWfwrkTaWCKtRB263ye
I0PZwvIh7MlZA2R8VvQaoo7X7J352j4EW0C/CxyWc4NlJXu+LmlXf6jr9Dm+ST1sT4pjdStWOYL4
YrRMLLY436wpl+lZAuJf25QrGczJ8cbEboAooLuxSRZLPnCIZCw3eIG8/lZ5/R3VAoxFjfHz3uLK
uDarItvnvSY78tzMwrIeX8zifmTOazSnYYkGBOCmvxNFSu4efZQ8Y6sDGFfuALvn2kUHHNjbBp6A
9T6SBtpF1sX04tHXUZtu4jwK+pmKgr6htOISIMI3VL2YIyb11sMpB1T7anEGkMqs8cvVNShXdhfn
i1Tq4s74tvlf/66BFD8W9F8saKNyGwtekJ02Y5PiywK8tB8Ifm3x6RHleLw+nt5hVvlz8nNJkvLG
orNGLJiJc87eSbmH4gUX1iNfqQR9YsSSKER1G3nJ3Uz1IehFrDISuOPMzJxqmCM0FT9NYMFHgkjr
qWjiGet0elyVc4e2FjIOdAFJNlINBx/E76AIWi9Pnis1P5nsA8N4Xd0OE/WhYdryi2pEeOHBmdIf
PV6LGXkfceOdzZs8fo5YqsyoDVA5iztRBiFz6/rgc2Xa2kvD5p4NA+/rvUSWji3FEE33phqNj6+Q
r8kDN8LxdqasjXg+5wu5XgFgE6jYFxlbX2Kbb6ZQe5eWVA21217I9iVZZvYjMoZotg6dJaNcT9de
IvjV5shCmSJzQao64APeXhJIwJoBHIcIIII6WeNdjHd3Z2coGEp5+fFcVl7MgIMV0PZwu4ZoJQZg
TjxIypFW9cryDhdiEy2eaARwS1NLavGbVn8EP086lZL8CRHsQGmldzKv5qcA543hqy+cfsgRV60X
TC3MKQbaPVLZSCX14JzlO9dAcNl0A88Iz/IchhrS0liPCcwDdj3qTF+Qo/LcrbcUO9OGia3M3vJk
+9RP9Reti/KnZnluw6rfjJBUs+XDkOqiSfdK3VRcgogP/LP04KluXenDTX83C2WUi5gdEi4J8qg2
6jk6vXgUN3B04tFqwyS1thgegJRFL+HHHfZoFJUAjV5F5y8S89QemTPXY27VcmtSFOfUj6tKxnj4
3gq/lMTVa8xr8aAE/PUFK9tAFbazaUlQmbtqR0AnEx9TNGbjR2xo4s/HXTUKxu7NChRgKoDo/mSe
PU1tYVzMBzLrX3JL6lMyU3P9h2gFNuyUPpe+0UMLh5+Ju6fcroMedGZL6TxZptibnuPBb/LTwdnE
/LxAngOhh0d92b8hcpm2m6Ax1ThVBNn2boioFgwRjzKvyY+sE79jG1rC0fmvQzrl6q6bZpl52jhp
B/u6LuJ1bOalfTvGaANMuqjGjfvl4afY+TA4FU128BjQB43486er06lzFq3OwccH/t3ayp/4sJCW
qmp6mcldas27cqOtS1IXgUYABbbv2GcQfJCMjsrzn+jiaaPh9oExrKZeskiu1eDwltgKEfM2gLTd
LTVj/6EKMyWPBsbaMIRgfQiKF2mPFIcVToncuRS6VOXfZbuRO3sgw2FdNGExZWNotO5ibUm1FCWO
5WpOEK2VUR3F0Ma6/9WUP56M6bRXZtjDUb4o/elIYvQd3b2MUDeQ2u5GsiiL+PYruDY4z+fAfc17
23Xo9lx871ViigyKtGxbFW62tUShHslWCO6l9lvSAc226ab5SSr3h9aOPVefJ1NJIyeeTn+9qwXo
BGroOCgEVXGK7P5ZQkXwbM/EyrZ5vgL+ZbHQnUFgmQ/gBvuSW/6HMMAqiXX6pv4pB9F+aqwfcCZe
WJV6z60ePlmbMC7+qgQ7YGkX/aoMsMAVTpnlU/ne78mVP/JoebIwcZ60nRKxkyH2WviXKdkxq5Fy
YVF09Mjvj+CfUpd2qui6dCiQ8a34InolmKUeEgqhLGuQhaauBN5EluLvVxWsXyw2qREKu7zr5YDC
xBlUkZY/60baDK6wBFUqRScAfOPZrCryKjgiQdadVWYkn44unqbJR4sGpuR85ASZtO83rBqg5QOp
yH4YT9/UC/UEaAfsZMDaFv+tIIGNZhnvnneP9lZHtaPIKzP5XvbW/x4p9f5IDE3trgmT/THezrjI
qnYgobjMe++lkR0s9e5uTAhUGaAoRVdojIK7LNaJXEYP6jvpY0SUKbIo53DtdAGG5OQnB1M/AjbY
ikbdrlXoYkrAAQeVyPq/Nck/i1OecegwuVyDrN30MtItXZGyTy8nQRIpPJrmOiimTlNt/2QSDtDw
oSnUrEmqbtPPYDxxT/o1RcbvYYoHrIw1axVppJpNUD1NvGfJF4p00hjXjW5vxw01wd9ygbMIeke1
HcJqaG4pg6P6RDTXOEFunR/iYSaP9adUjLzODMHyUPTMWBIOIaTh3zLVdn690eiF5VUU2MRG9qfM
1kpjhOKdddSk4TxtOXFrCEI4f61F8bIzhmWY3r84zvNSZw4Jn0W96lYwqNk2u7ohfHFcvShRTRFX
9nwyALdNx2sb8YKs3QHCBiRjrgtz7S+OVYuT6Z+JF/sFCqCKYi+fSBX2DXUioXEbT+mFA4AuMLWv
h05gLFIEHilCddwTrkEo3CoDG35f2hAJgj44ThP5KJ6b3bwG/ncujweWucH2q2hua+xkrvPyeDzX
ggCzmKZz/x5XqCJav2ulNueNDJDFs4OuLm2+4OSrh8DkIi3Xgng/J7xR8wF3UkqZV+kZ+R6ysWkL
xKtDhvP2M4ZW6iX95tOR8Hk4lcsbJc2/BgRD6o5Q25S4814nZyTheFdSzRDDwp1daeXZw4n8eRyk
zquXLh//amAvxuuxxidI9Vxblu4leRMgXOM8ELwR0KF+a+NRsBeznVembcXC/RgR+eqlvZC+tz/b
KmGiFZeERnd73/q0ll69/iZMIEmPh6M2htlt9J0DoZRh4Ycf2HBB+YrnoiXzdAWui+74V6LnxSpm
DKwNrm79j4ZJ8oWd0ficApusnzPb0J9AXlOGqoa02EmiqZGBTZ3oSJ6eRCzi+1s1/nAt7z9EYJTw
ZopqpU+GXo1CtUyc2My7CybK1jSjZnOjjTOERcFHzpB8dqUXkR8wCDTZdZS3YNGq5xhzhKuqgSyR
zZwGtfaaJVQB/xhI+0yTUT5PmAzT/J9nT9PgCk/05jU4I7bZwAD9rxz1p/NybvLGV5TatcOsmXKU
NvzwP06KqIlnTk0dNPNM2JS6Sy4awtdcgtL4y69zc16tNBURiC/GbVDIWFqCaf97sapPM1TyRrLF
SsLqN25wOadqq3VSUzQ5tA+MN4GXKmTeiJjVziXmUF5eJRo+rtA7DDq04tnxV4N2Uy6EbHg/R6lb
2aTZ4yppYBjEGEK3aZJVz+p20gpfLjXVeVuCNLMMVTYgoxEGZY5MqYsqvk5LWl1lXIp4eX68Rtev
P+eev/+Cf0p+5R8AeaiiM1Cd4HzImwxPZuYYpc4/XXh3OtywC0oUWdOHeRjCXTGa13W0OteAOnYX
NOFoSu7quUtSSEGVmwg2FeGrRa2TjzkZSJU6FVqPnCUldPm8uDBMGcrFwvyuzz4r1as3X8j9tJWQ
IVGNnmLW5SakzOn9Bkq2VCdy16v7m6ZwVtiuenGES0u4+oDO+JHZzcveWp1KT/PiRwkv/cDBl5KD
ZKgpmc9tcUFJyEEMdhcKQHtj8jJpB53u3A/fdz3N57qVgpzlXSQeRnIpeOC6gYyePtMGrPUOX9lv
DgCAfyHrIU+6FTBSSX1K/AqliRo78QuHY72WRctvVngn0GqZ6K+LrpKE8XKVZYlETlmD4XW09cD3
ltRgVT6xG+zf1iJBI6W19V0faJn3akA1PlC9mpoHTb5INmBSIUDahSCwpYtyCvEFtgZ6Ugf+5X0w
JTtYYLNKNAQ07niLUjf31CnVt2KqM2TuagVoQfKj8ruVjLw0JczM0REr8vWRuQVwdpO8/SEDUvH6
wOaDSDjR25YQ5D8Ghg6SQcZWuxRdjbkhvNUykAwc5F471QsDHhvqW8PMXQ9wa9Kgh+zQXtauiKuY
+zCYgY4Dt2yMPQTHjJO1kjTZtjynhEhrcpA3Lt/N5lQjI/nCJd9LX670jWw9c6gYTXdVOLkY9e/z
CU5YGrVMg6mLJsp7ucRxdzfJSP0qz1YhrprcaeL3ybvO3rtrmrQi+mifPRFbMiiHQZC/s559KyMv
xOAzkAfMbbeb1ItxCo+c3gLAw0bVY33QeGY1XNUNng5jeso+aBiNycn766OGaiYi0/xVSJeuOtM9
I4BYvZyvXxqScnzbw0KwZ2CAOwTUcGEtHUkoTpCi1d2s+NeHRMhH2gKkSLih0qCVKFndLP62AasT
QBZTneFyV2aDDm+708FK40rcVWWcG66l+b+RhW2vn4kP/k5rbG5cf0UgA7ADvh2E/XP5geTiaUQ8
2z/Mfp5WKDd2iQq2bL5GDzYK8A692xKdpj0WB7/luC01xMsZJJEEZ6i2+I4HoyqD2BL31O8OG8QZ
rPls8Az9j+s+cvgF6YydjeETYgi4hsPPinEqiNwjOc4u3C27WyAACHTSupSERXINR0KXsm3/qZmW
VASdx9MUt5AbQfemnOjrxe+aQ6g07l+a3wmAbc3UZxWKhQZKdjHZIgKnAwm9WvQ4wX8LstNPyi6n
AhaxdLDLT5G3rE60S5mfqoaMqG0Pr5Ni6mF2jrtJYrzjLrr0kX5Y6VzES9p04hnLps5SfIgC5vrY
Yv6USTReSbhvadEmRruZu+4Yh8dOQK48L70hm9OKXL/mAfahuiluLINzAGCM3DloFi9s6iW5D1iw
jlLreBAyrioJcPTTTLiWVj80dvvgVUWnFlHzprUyyp2ECX+knBpY55eo2pSenvPBXxir1n9rfNdp
eOFZvXvu9NTqCkR0R+KuPxKRWIZKs+gpGeiSujbc4RMr/Tz92MLdIkc0/4loibiA+wxYuXZeEkf4
XrHxk3ef8MJ1Sdx9iRwrVx37bNFjLAsBo33n3NoucMs4tqTTH36Vc7Ri16lWY7YhjA8mKbUyNEpN
HxcPKboGqItIHIGuP4dgmLcPUjZg/hPOe3KfpyeixJBKHjmXHZ7mV9veP8rEnJtIsM2apRTJYIM+
H3HPYDnCuct0oymyMqB9xRVB3kHvKF9xr+fb8M5WV4gwyt+RtR6wXNfuAsEf91ARiiv+RBw1kg3N
ZdWLUiguheEjhMpD+vPoY6cbNccM/82ywuu9CUvJuZZW0/Z3S4jmXOQRil8Jkl3buRGnmAx9/9B8
DcwsJrZNl/IV9y3BtRIf+YM8+jtFtSiZv9gUUzxUcen8iUmviKoJzXPMn1VSG1Wny00SL89CmNOR
vm//EFCxiyDZ0tpqUwZxRnuZ/hXUUn7HZcu0oN3o5Fygdj6XPY8FiDgaSI+69mWSYzvUTw79NWkX
MESYNQfSwG06bv1Abou90ki5EpBJ4iFF6XxhIPp9yK5XUIw3ySg2l9JGvKzlTMM/AfGiY5X6KoTQ
CR4ahF8vhv9XeIj92zC+SDCsKeYH6QKQ+VJSVeEgxVtifd5z+4UyooZD+WQX+wgVNWFHAw5ekH58
eSFHhewRajsy5HRxpTb/AxGnjNfhsM9rNnCIVTwOxbmMkBvdWp3cd9o6aoJF/8EPg7ZtivitnFzp
T2OFWnuuH7El/mN+q5gpPPyoi8VuQbNk/u1TaHUSYh15uLEu8aklG5nc/OdKzj1jHa3n6jI+jzEI
4EvZQ6y11x3rgAJEp20FcHXABhcy/wntWZ9CHkkX0CH6Cf177ciaIGRKhsFxF+nH8lNAA8hqlomK
7izxOwQXkJA8sNJFdojTGJAjtpflC8bYqjDlxVLqw5QFiEUqFQQGJmseQsnLZOsFTbkRbOL4X4GW
ba3M6zuwEgcJ1Mz8WJL4vwCnHGnOc9pnaSM/cnwmX7R8vjStC5OWfAxAWin5MP4sEGtdi+QuS7eT
vgYgJnG0wYof4DQa5YyRV28e3VmGIV7dG7JidoA9zrv5iEOuRKegByZLkFMNSgxKMMhI/psLL6Ww
ODc9fcfq0jgpnW3dC0tqVGJ666NARz94oMVwFNRBmWtztvcEFYKjY0jV/Tp8Zj6v6VdABAj3/IwT
cbSa+HbjQoYfJr8vUxwwcHwAGwvyy0M2vkErEWDLCFbLyWu5pwfvQt7FRb1cXsIqIDlEzXwBLICw
8nqUoC2vpWPIlD9jG68Yy2/Uhd8r/QvK6lRhUD41Nlz8dIXpndlVDQow77XuRmlo6i5WkDZFi66W
T2UmpByJGhV42dxv7NuKrObdBguSQ/j1WT7BwgD8eNHVV5pHMkHv38pkiw7es/DZXzqnJqoHeCS1
at4uzbrFxBkgucdK0qAts77rtYEX3mkiW90oyhOddOHLW3RkLr4Z7X56+gTGa7rKLEToLxzNIDX3
4a/cXNO6nZFCkR027FzGXAS0BCMqGKMN3vOPxX/awoMY10Yq8YQGvjoNczsMnIFrnHuoncCpZP+s
gqSJgsviXNWVLOW5ftmadJ025op73CYbQ9G6cjU1Q29oEoJCXnR5N0rzkaA7P/BsYNtJQpGDaNct
4maK3cUeVKx9nZGKRKyqpjNvw1LZuqvlSO50ZZ9auWw8w3QrfCXtcX9MD8ZvRrJ3sZr20arSE6n5
/8DG5XulfZyRANgxEXXoeUudzKOYoBGF2w6GJk/RVeiB+GcBAzlZIjHxg/voKl1xCFDotQNsyTnP
SidVY05lyvTjAd2TeaSxc5NdLLQthxG1/B8Fq+fQjXy6b3j9GkbjiEgQmZtwnQQe5UgfCiWRtCcj
2l8vRXnWWo+w/OrnvFnUu7O1dc4/eiViRb//K63FrE++DepPYu47v1cZan/Cd0CfhpcGSqahypdX
W8ruXe8QA75wIaPzuzA9aZjUpRKjW7hXdU4kdAI4PGqk/dWu3893Oq2oWYGudg7l00PpSR/qZ+fM
lKtXjmAuEysPXsTaen+7FhqCWujCtY/98WfnmBlZWtzqpp0Isp487+u9Fwty+CHEI98ChHlacG/l
IpiU2iOCqT10jwmwwfCNd1uuM93mxoYbCJuIuBCkXskh8P4+g4eF4aXLHqXf0o2OiubLI4caB99q
p10nPv9AmHw8hQBd+dCFFODQasmqpDfxmch5XkgLGdafVEt5ug8ZDCr+aFh4KynmumHjcpgolqfV
K3vzjElQU+BD1TknJjIHcByHrxW8dOz5DN8OfMx7rUzNg9u1zmyEfHJ2TPNhX7KGBnLYCzMUJ0qg
R7nC1BXUeqXPKPezSGmKL/dGi+hq1Btg+C7FRGAr79OloK6lZn8PRIpVQOjSCYcuOYnpn2EiJypM
llb0kz6lDSRm7l6oQ8eL5n3E/6t/c3NTUz88Pq4+dIU3h8jovRgoSuADOfwGZC7igCjWrw4rIe1Z
xRRuoq3b9nimre2OAEVj11+SlX4iyFxkdkyevSJCIp29PW2bieG40bbCtNQHgHE5OAAMLDFpAnoS
nbxDGP3pXRMymT72OcwPEiwGin0d388xhKYpfbEftmx4Taif9rtZG+wI3DJ2qccfYNLnyC2Vg9Lt
URETwej2qRr1q0OII3rRbkPx1T4Gifewo75CtG/SbJBD3aCKLRPGM2oheIs8EBYAlgLOTRwB+XNA
9RDqw6gNxm8gcCWbPzgmFYs28hE11Ckfl4D453dENpeinHkbwO24GWvRNRYy3oA5jnvKaiaa5AuH
40AXvGJ77J3h48yE947PJpNOZeaLagng+t8BuU02Riba/LdACpV6vBej1EUShNuFNNfG9lWKeByl
45F1RkV6ClLsH7PUcIwwwEiYmhRusM6QgueAyUXDmT31Tw9YsG4XctPF6D7EFAaqmBt8UbHL/J/B
zMtBrt/QqOzOYmvAtrvQcdKmEpWyTMJvrkVoHTYj6KlrUn9XD1A8b2aHJsf1/7+rCK1+/IiQ3/gt
gOHNZfW8n2SCicMcteijAtmO45rpSIVaERFmZI1FtGTdJQtkjMy3JpdGbKUQubLWyTh4NHT03Tq5
1DKv8pGaEEZOdnQfe1j19ScgL92Mz+TWqmybOltqXXwwGxXJtMHbyFIyAnaWua6HeEs+K1Yos+gz
8d+ippvsOLVwOtR7tUEcug5oiq3Ap9otuHLTGhjcdzRrbrk5RqhnX7ah9d1fT5wesrslPPWg9kad
GH2lZM1w+0t4kyHFfMms/p6SOZ9LmyNoQVSRmgXStZvPv3hwVmhCBeBtO5BPiHwKI+f5NE5aJOOo
08isx7A+MtIpKPNrhqqdeJ5E0ETVQLoGzwa42OXrsE4qJQxCaMNyOgke7I6A5S6vfyxRzGkrdI3J
/NyGLymdzpWElQOXSnJSbRxjtEp6wzK6yxo4BX2kOys9FJwRSJtnEQLxhBvuyYGPKFByN1NQ2nue
KmhWWvH236yLl0gNsexv6HdIfGRCUFq9dXlY2cEcEwHqON7z68wAzNLdNWjg/4CsgTc3vZDFUsEm
qtARZrXqgEr2CzafNhhanHpbGkF3RORyZdYW7wcnd902t+RPjuZQr5TBoVBf9hMUAc8kkh3biUVu
KF6TI33Q2ZS5FcuV/+XKmo5i3uUAPMOEFO64QM5vgTufzFyQIhAtZilynplgZxqbe2XAiutf5kaY
ZbJvfi8fIkPKq/I6iMzsWReqSTps1NvOpeOzWtxITx/x2TrxX4OLNCfho+AJCINXAz9FKUVjj4Xd
fpa5qPKG/hhnI2o7geM6SNoXlTr/DTBmljGLtJ9sYEk/5HifAFlKZHp0nEdIys8jdNTPxZBUP7z8
PlvDoAPc8DPSKcCYBHNdiLausu96RvVeTh1IIZ3qiiPYC8+VGcBkR7bnqWdsZocNGkllQyPWYVCz
wwbJJeafvBJQ1U7u05LtoMy4KuLKIytryFUdoaQ56ctBuqURuUs5zRTXOQ5SteFs464g+trNqGrk
E8VxTT+I7dGxge0J7uKaVXxgzaHfx6Ym5Fc1RbVjTBQrI2ucBU9Dp8g+jIGN7Qg8u3do1q64Oc2h
rMh9ghDLzQKZdWMsLmupobub9b+KLaVbYVTY4INMQchm4TtqQrE0iSxJa7+1CxuST01CyPKsjrkN
alHIMQpX46Lavd3M7fBmwx2JSA2XTbRphv3PKDYO4hlS2lvbYTJ/yFaZS3QZE58Ina6yXkEDjM2O
0RDEfiB3AYFGRg5HzGvUn38bxARG6MZcevsyyOQVRD3WhRZDTTZ5FsSu4FScRhHM+mB+2MR7VJ1D
a59hHH8XjOuxZgIEwMd5pp5mGNDvWjHWI2YXEQL8AZI9upibokKWB+iKdvOIIZxsasF0eocSgrSg
n4llJvsVgvTU5BqXbbE+j0YgPBW7bnG2GJAl3dRoU9gZS/vLSddFe71GZGl7FlJEDDMb1B4d4eW3
1jg0VG0qJyhc68vrZKxDKqzzgvYGu+1kmdUaRkb9g9hej5eLi/W2bXIe/tW5VlvuqcAKYExH1D5u
NPQcHgkiK1APVxZPat55Nq+VsBXQuIDOKC7+hSUC8yHYIXodplpHm2M9gNaLtdblLALUEYpG7yBG
JW+Nk4mD46jti7+Q4NXC6EXggj320XbwFDssdR++xqbiKzQr4rZddGbMEP9hOauTt2j3QbowVnV5
jsb8GHfZMOZ6akPyIr7vocRooRim2OZZI+j5og7xF/hvvfIXKj5psED06TYatZktDzOPzF6ZxUzp
1aK2HylymalAGPn6m3qZwCG2Hc9QssTR6cT6bp6XFy2K04bEB9qGz0o0xZ80PlQZBHEWfvYl5h8J
nWI4QBRKuQUI3BjaVtK2/r/BO3WAckPDAYDv+Nt7Gvpru2dUxAqaDXbx5NPx17C6Oj/yaMTnt1OL
JBlGoISSRO7S2TS9I2sPTel529PjY9shFeh2OWLKIasMv+1BECYftFcxTXfiPv4VMss7+ewBPaV4
iYKQpGmme5iRfBJVwlXw3EIo+bx9RkpaVW2cJnhFAGtyFrI5cQumzybsYd52jBhrm7SuK3agBkE+
io/FzUvC+vqS/kGJfPIEbOPjIYc3jgz/HtX7JVsqVoMbaEKzOlBzL6T1S99jXIhFzGhpTmlGwl3y
5OwehCnyvycEGep+m6vOEOq88PmMGQMLdfcbJP34RwzUIczoKgi/WRSYiGP3dwFUC4QwT6gHjLSF
p8YpOkQsVT44ze5W2Tgf2IJtup132QhWq1bTimYm3ebGQ++nXnNNRpdsTDpU8Vb7vE9QYhR02d6G
J5yU/JR5Q8TXLVviKsCLHSAXnyJvComw4Xfha0qZjNpXMr5h64YnCpQ6lMo9hFF3UWVmmoufMFmE
RPkKioTRmee4fvnjcReZESKQXM222l3uvWDvF2l+HDsdqr7N1lc5qq2Oh6NKDTuky79CwSdCeXCj
592r9/YKw8+nVn5ViTllg7awm33y5yG0hMLHL4v5n52vx6qI5Gl334NA0GNBJzFN4HwwIG6mGXlP
zIf5WKhtDJRBZzwTIn4xWmbyYP+YMamn7VfdTTo9ZWUkRvS+pMkuWHKCjz+HjeamDHZtKgWm2rBb
3iAxrWbIEXUCg+6sTWfMVcmi9tInSeCnHKmf8i5eFE8FUUTt3UmTN7FmKeuL2ZAVh0D21Z5ATqeA
UloeHmYnzSCsUJXX4BVMACN95pxLfIsTnz1uSUhAq7zJ9CDVxF1kTW0BrlG/XIYvJL/nHvVefBld
l4duKbo408Mqif0U+buqd7fh/v6+ycx4ST9B1uP/qaleeMG7GHp2y6eQ5fjE6ZyiqeKQrqBPmxYn
SOskLUSdWmFkIf4cerq9KfNblPR3avFExUO47Qwm/aRPiMaSOMNFi0JkzGiB8wkRFSSO1yQrRkX2
kEt9lDRZbt0AqYqqy0Ln8TDVTx2OqnqWEWvGw7TJ7ex9ECX2p5Cz2lOhSl1uFxbjqUp3/V87eX+O
MHQ3bX89IujG8MjJfyBUx6MpyjL8QBPX8TxQNfSaDD1ukiuD8P/LOcZZcI+Mk1vh7Bv4i3n/EwRu
K9NMGRgAhdej4RmfSvfzG3B5nupMt1hCUXLZrkh75os243KWxpszqoO7m5nFs6v+45hW/B2JwQaS
BL0UtKkedp2BJLLOxKmP9rnbgSq+q7nqHUb9uWzdcDF8qukbfOARU9oZ9Ss8zr48X2RuilS/jUJm
XufQfTZ7Y3Y4XjDIYDy3ItEQI2TlgW8PqIr+wXwUPIrmS39M2xkFl4buI0VxAYhqjIB0coviAqET
p+gcJ2TUQh/knukT3TtTGMFm9gn3y2E5IPL+i8Y2aj9NnhtOGVj/3/CHHHNAYmFZn6t+otba30ni
SoqY9NWGvlGDWthaOF16fyTZ3oJGtyalGHNiraOQgrNtBdegY1Kc4BpYtPPMqCNxOXpxru4sRLCo
uQGfQkxu6JpjmDvqxQgZHQ7ktDh02ZtFFt7QtwqhVPf7SN1P9084H5Gg4oWxq/pIy1C6YX7SNtjT
k8gYnDfLvxKWPltwt97FBmF/RPEYO2qRnjPsxflQbNv6teY66m8JKTl+hIyspnYNbc7psFPYrG8o
iOAYW1q7nmVrkU23mKxLl36BRsLIK9h3i1F8mvFu//y0TFy2dzo2JzURWlqOfsWvPMf56piDwj1c
2GUvhba7Z/0Oe3TroATCOdGh4Am3yz2fXCkzw4TegnHcgMMEM+xCICr9aGIy/nNwb8qmW9Rsi+Iz
Av7V7+EGtP6D0KLJXHKWlpmzm1q45DalD6jL5fTAaZF+NAYUUrUD+tCdAablrQt0p8MN+6biV+SB
5AGXEUUUa9RXRAgC8dvEbGy9g2lo4GfMsJKmKawBHoWGWR+uRq+GsATQ17pNyjH0Mk1j33aiQjn5
HoFR3ogKbbMBWFELePwuHAGtBuLtliSQs0e+yHPIgFL7mXC9z3Y7b6FE5dhBMw/d16K7HTLcYKrP
UTVC1g+rpFkcdU5z0f39IQeVv7JpRbuPtD9AGUC2i8E8OQs1VRYv8aaJoccRg8Lv2SLtC3ZrqBvQ
4KN4NXm1Gz9q02fXYOXlx4ALVRIwqCYm8nXEGUg9FEMiRrU7iBhDNtnlP6HMzprjxAjwjFy43Tw6
vq01Vj/H/Nk0hZIlrjHWMyclnrQ1E5dfN/0Lv9JGJNEuT2EQnto5KUK3hsOZGMaaVZASGrK++6+j
s22h4PNsUfQ758SAoCSa5kAK4tSlC5vWG1mKaFo/7PsE2udul+ZmX1RyAEsAEhgmx+a/9oQ9XB6R
uaqiW7Jo6RiUqPC2f4jNlhdLwUqjmx0rI4Q8ZW/Fs1bu7TmjILPsaO1sjpKxe7IWXmIeu8OKbUZY
IY+EWvqOOlbx3XSn3F6QQG4wBn7K9UHVzvxtGfnL66Gsvr9qAtp1HQQMIJjb7Vlj6Kgnl/uUW8LI
bFv4PW0/9gS7m9FkryZ9LuK4sX9Y5ZJzCRb9WUFysJERwEf6WHdYtV/BzbG+HF9+xZY3EOYjo5Cw
Ll1R0ZNPLm2n2Hnmi+LdcJZz69aDrDC1mZheFhmtq2480iRlbePopeec2DlWoyWQ/xiEY1gW1E0Q
XA4tBcp/a28U2itncrimKZhDZUQ3IHxp5n0gv9/7a49Bl7wg1ZXX6VzzM5P5d6IusPEel0/s+ASj
bKsKxrFRYpWZXaGO7EpZl+H2aboAt5s62Onfe6oGtPNJ2JkxVqHxIyxFde+kcAo59TS6JGzLaTVc
Obn+VZDS5kejs20VyDLhTHJ34CzatM60HduWsfcSyF4D5paZ1kvRzZJpo4zpIUgxAQ2+mju1TSgQ
Gn5kud/8r+uVqq6Yvx1hqBf68oEI2Py+mo0t36UEeZ6pMuyLH4YjbzjTRfvqoUr2J6q7/f5eSR74
1CqWh8/d8omnudqzm5IXqt9jN6i7cAJkrpdga7m9Wr4aGEOw8LATjJV0EwjtUB5YRi07jqggEQF3
MQ1p8IhJouy1tO+ePpvIVX/+ioZ/vpuxUNjKsVnJpk/uqG1XL2CeLKR+1GNXWKTvvbewrs3lIdWg
RLkDebcH5f8KEkHJimlmJDf8oUbIjlt5RfBFcpJDBN+j2kOgCfWVCyFR5ruy42gSiC1N7B03jd+y
KSa1oHVMaGJOwPZ7Buy4EFY0IYyYhQ0jit61pkXsEzcPvO3L1RSRjkEPwPDd1HMa+ZNl0r+inOqq
uUy7od8iOpEuL2EHW44Fn7uquP4Aji28ze+eDc+mOQqnD7Tc9A6ptBkweUwJRHfUdeUM0wij3pQ7
Gu28Nrx0NtU3eLHooK8TE2Wel5F3khp02yFtTqaYmsIdofZwzzl6yKk1G70GSPsMrtX/aLEs+pJQ
fnd4WjlRkc8cxoHmTG7bgmK4OyKtYVyCxsjL9LU+aYAnuO6AeP8u3W049PdXa5ZnsgYixtsCbcEF
kTRr5jfRoua0t4It3W8HcHx0WFDIvaQE0V7y7TjmO5uquA5W7/zrQAfP5hp8hcVS789GQEW9ukyU
5J9l2h+iDV8c/JEPIAylC0ijKnOiMylX5bA/FgyDE8vI+xSzNITYO6YDrxMazgKBR+j0oH3eT+nJ
xPmTDLrAsUIhkTx8D8VFbEfkHGFY15aDP9DQysfC7D1GFj3/ntMq3QQx/tEEXKPJAsDcVbAccMhZ
WivO7MDtReD/GnfJIeYjFSh1d99w1wiLHXCuCn0JUEQY49OIFdujpjtxR6kY4f55NrWhQUqRty4G
LF1a29ASPGdLvi+rJMp6ZcgpYdC7vpVzjRKrRFW5qe+EuD6Jy8LP9jPNhvlidWQSO2tD5lmW2qvD
j3vhdm4rCdxfF33CKe5mot0oKpeRtB8BePCNLPIf0GJcDyAf+NPMBylMLOqwrvEKhpz7Wjdg2/mn
/gJ8BjqcdUKPJMeLXpWZQbJOqtHkJdhtsCinvnUC00/LvbIkTPlQMCb0sQINM+ptVIDkw54EqolF
0BblGdpUw6wzY/pEek+D3JNf2HUWe2q9p62DhmbetqUYpPQjMZJY5yYi2mUluaSL7MZ5tjDj8SpY
IZ6m0pIBrcwwEotaEAsT9VG4THThBi+5dK05FAGleq5QXI6042FpA1UtnWTWFcOEZKxn8Dgd4kaP
jANR+rIXFkVD2Nd6rI2E8bfe6sQdddkccwkTg/0IE+3snmKrHB59wtvGIxmxhNx5eMz0gsfCvN2j
zyNKyWOQrj3xDxOB9f3JPD6qbM2u456Q43gMIrxuULIdjFgHSlHpvcSNlquzzy1oNrHNKDoc3YL8
ijXqwRQVmw+hr5QFvOfez8mFwGij6bBp6fpYVOB5qMqPf+NSN3Qcpb1aKono6j2Sdil/I4U/d8Dt
9g4J9/+SCgsjL/P5kAmzsZNytqVYXePRHp7dK/oasvFPebJ+A8JWauM2UvjIgibjZit5gzIPdQwI
tceQsrdmShPSHIFsTVcrw6L51gJSr4S/Fsj2PXsI1kUyesFrNTWAy3/YqlRMUePjIUQ8RNTg361v
ngttDikd507vQIYi8ZE+Sf9u61uJ26Rt/VxoN4RLZCYWOYHy/4Gs/bvIH0oZ4Mdjtfsdk6JT7H7L
sjEUr88xVh66xv2dkiQa2tUucq0zCcnFKz2tmg6f2KN3RJtOw6OhDAFGqtCii1MdhKsKNM02HodP
xiTvpvAkF5aTdVFl9tssAhVImwQd0W3IUnQcxvPnNKUrawV59PZUb/fuMlahFtT9Raee64djzqxr
qXrkRvoejfxR8LJyCP2+SgSUpQrKYMqQKYg5SH4QoO3ZHEFQwC753IOimpvQAgEKlxi7/K6snm5R
XB931R966g1WdNxaHLNWf/xPFDHGQcCTHvnT4ZEocGDOC5fMfgp9Xjas8LqGikPrjXRm+/XBepz4
G1gppZ1TRcjnsHnnM16disY+j3dyVFQxgGDi3rz4Idd6+MLWb9mrHxL9q92qw3pnq2TeQkoc10Ji
f6HlSfCzNexuoqG+8gFcXKnRqOJPYP8DRnCGSSFX87+KQ/uwvtarsCifF4649qbaDPJspMDfgN7I
uIlFHS4095vgVSDmeAmlM1tjUUS5wn1KPl2h3y7m58QIprWVeD1T74djAFmhKPYiSEoWpENI8RGy
kXykSDOAWlNiRXuQQIR/bZfpBfVemk9Qtzkvyz7ZyG0GJtlBcO7+fdeVvBZoB/FhONLkYyMe61+f
CjWbXmfugzMtBJj8iCJ53ytIA164ExCDokzpnpzToTx/7I+ia0xVrdvtph/NkfaA2SIzAPaOPdqP
gQBgBbQxSWngAAb45Z+tv0ZjmBwYrsMlfEZ3gJT4fRli96DlD80hYI60uJxFS5DE50H/7F2lZljo
/8mp1CPDaws2ZZq+Z/Gli2p3cKvZj69ur+BA54BB4kuOTQpir2RTrUprSHeXagoA5m6oyXYHlUkw
6RQLEJI2TS4lo9n1fD2X0J0s2RfJ0t1s8LGGBjrhbsiXko6kageAJDnbBRbD72qob1OCBVXp1I+6
Xs4pjkK6JK02jTSovwgVigx6AQNtdJS8qtq67LHKIKvRLMZ2a2QHI/jt1Uj7rzQZy62H52TuW+Oc
4tuG4Deb6LYzKFknA1on8zhRljW1OarZiCgC1m6Tmm21stduc3PMSTfFf7LRhoEIrkUP4eV/oWLV
acyM4l8EAkk6GJgwLMqPgeK+iCLqa4L/nYeUUfWzi+2kA5zOtCnruRhQu65vPGwlHzi+CMfXgVX1
/OI1s5FPpNG1C9Lg7Ot85nWvygHyJSDJAexTbE0Cy/X/UvBEPbILL/yb0zJ1cilZ+NDhDyTc7Fh0
MnI8vJg8yDjgR+r7k1dGXwbeBPKIrW20/eTkBxQBWCDMzSuBGUr5sw3zqniyZuXavgnl0Rcnx/sv
6WonplU6JXpanKzuMTOiMwdE9ommbSGc3kuDK+mwAlGCDFqhXu6I/Er/KQwXjLMftTuTKLgh0ajI
XnG9pxIwsQqhb/QIAL0BX9h/6SBnKX/VymwmWRly59cvnKneZeFE/u0QLDAvkC25jHOdLu/PNXWc
Bp3MLr5gkS8/YW1q5Dyav7B87xS/oU4FxebKgNeLSRCKaxYD0O1eWpWVMAQglxK3VQGDAPGv7tm/
KPv6aVCDJkOgWmb2MHxIMdJQxWc8aXKVWanOZknw4cKUDBBOqSA80FJZauFimbvQhCT/lIx6s0d0
uIGk77op5k7Tp+Xt3PhlrpVOeSoFT0/OA9WOwbwbq+kdFmy3y/AcfmoaN/bjwmaF8gQ63VL1wrH2
8w0UMi8lDepjjHzd6u3dsgCvRyYcfQsW1iwqztoTTu8Q522egpdcFoOIZacdA6ZtKvUrymP6qPpe
bNEFBR4TI9znfa5TPy3zcp0jMhqojLNU8vJzYrGXVOSwUfVVdtIJlwlXvJvRfBCrHPuM9gVu3WpA
gISeoOEg7aFrjBuqy0xy6GZdcSG66oXinDsHmHrTLQiXJrWSVZzuDW/TFiPCrArfohpXB5i5EQug
TdWUZfwUeEqE0msyQcBb7Uh/jtiKF9mfRnEZfMAUdkF8Bym3MaIPmpzGxfTMbPi/Ljn7Xy7iulQV
1GplZHdo+0oWWsEGiRvAW03UP9fDzca9qkDrG65a+a8fPLWYDZF8uE7M2Chca+9zjTh308yZ8lKe
OJmWWvBKfvx5k8N/6C+cuwFPk2XJGu6IGFQvHeMXHHeIdqMwwxcJEJLtYJk0tq/dP0zXN+MkpTZE
KrGqR3ZKLk5kJ5mBGOJtZvCt3xjlP5+8mTAQUL1vW47pLxkM28/QgAeJCTNRgTq4qV91oVxyJOb/
uF2ZHk9GA/XTGG0wBmK8qu5ZKshe8Jlwjy1b92SR0E6VvoGlIg5c9orS2kpB5cNOElGVGp0+qbgN
G/FmSM/A76+VLKSC8L4Egr6XXyXgcWP8WI/aKs+oY13Au1DbA6kIstJ15JEaEsxqliG1V6JZrhpV
TTP2M4u6JgsfAszadUu7yDaQUPNrn5cmd4QaGAtBiZQI5qQIottk6wT6EUwhCFOl9OjjHUsCRcNZ
xDAPfqqj8zpdKzyyPQgeZJPBQlpopRFDDCOEE9WMmZ4uqpLkNWuKD9t3WtRpuhuyV1WzotkfVEl3
zwFPrCnrVs1d/Wr4T4Sfq38jk+WEKdk9gri2ND/yp6636gHzcrOpaYcG7a7AyByNP+yXTmqfLo5q
jLrJv0uJ2ko2OwlxL+1FMBsPNYTtx7BEk5XbjULrRiRHCpDHwNClE8n/bGH30452MXH/HqSO89Ui
TTyLp+BkpaOOslOLpJS1xpYgJYMT1IdIQGvhn6WBCUN1P1Vps6QKT2At4LONJdlwp50VVZBNi90x
mmGLkoK+wUhydPh89MVZ/hef5QgunNohy4V5QRv2qeImeG4oIU5qdb6vCGcaGAT5IQ6Cxs79WFI3
hQKOQz+eVAeinVnZuQm2DL1z8tay7leQLWx8YfUo0fzRpBdyzBepDHLZM1ejDvAev/Nciic07li7
9QsQIzhBXDhDJplrFpva1lSuESV/CQEEq3Cu4al93OmSGNlqKRqu0kcxKVB3WGueztLmS71fIhJz
sO870ECnGNIghf9EAcnzm/CqvnBidRPU4L0cE9RG8Akrg7/TUZOUe4oMDejqgIDfySTKa1PMyNTM
ys1P0OaYDoq338TNulhVH09AarlpL93VBW84appeace1BCW/cHRoYlxshDj7m02mWFKXn7M0gXux
oa4T6tBHZszd+nuRPkKVSNdMuZO3PHib5nwi5PTlFq8H5SzGKo1ySn9yKjV7IZkd62jnZz00sESP
UoSalZolwAgo7pXiXbUT3xr/JDvuenOdfofbuBJE/D2L4RYxpa+3OdE9+yOYUWFA7blStB79qqMH
/Ts5KIGKvXmIOff2mVx6tC8pTLCtmYruN4/Gqr97XKo8LE4Pb0LMjIvrV+dwvsz0PCW9uDjGzN1Z
wquZAth6lLLxhqJ/KLnWjTE2i1Vf+BFnr18VZGR7kR+UWFjFPo6UHaKw3eSUqAkuDUPkfiRKcq/8
4HN5qajaAodKcBg+MGeKG+HSaZw+9HSqHogAJw5x8vusN39Rr5S7OTdQhLPCiG4on088pwXGoqkA
G9XFFYsfvJa5QKqMCzcnvwW87UiR34qpN2M2ERe76wcElA6bEOw12wvwwuXd79Et8HkECb1UthJt
d4efkl3+tYEi0G/CEaah4jUXnB+smXTS1VB1DeJX80u70FBuHxb8NQt+oqjOFUDu54h3YnJWFHMl
lnVLsVN47cKGx3UNpMxTJullY/7CbxPWkfWidH9gxPUshusZ8uP+fI4wKNBeqnwvoJ7LBEUzwIG7
gmmUu4NFRs8YVIg5EpYEas7mdtVXtxirotPUKVsodK8o/m2j6YJa2rKYWFG9MISM6p2+C1n/yCBv
SFD7O9dWmSehsTr9WXTMb7dzIeRlV3KpiDQ4cK29IAElNraHZ6jhAmAOlLDVEqTWjHKmuhU0LbcX
gF1jchx1r6TPlFwlraAphIPyetxaJpjP0EikuCZj6ATWOGd7vKnbZxxWE+HBByBuOxo+VVQ6BWUG
0j/IrsFnLqyCnO/9pBZh162VwjJMDhqsjJpEJRT2bXzIci0zMniKQ1rsV1GTSJkBma0YtEq2Jh1q
fni0aTM0eErRpKPcuK1wgFTrqaODwqleJmvDe3mFZ9SruqzeQiYWwGpY7giTk97rloSekVxm2jFE
w3VHQP6PWUH8TiCmQbr4nLpL00aQ1H/9SGUEft/2NqKhi52+dZTowhiXK/IsZ04t6a5C9AV4hQhK
MBs8AK15kcd1FgtDCMVa7WwEt8UQgF1ug/lwuTgmnWPnbeUo399IafKMn5ZlTyhWREj4VdytAsEV
n+2RmIer6tv7Xox+D/BdJpLDnSmDutIoqrFOZykZj8q0VPU40M3uYFo7JEOY1nQB31oSsSbrVXOp
Kt5kpKuHcZX3wjr89iFrFNFRZQGrgSEOjwHMAmD5JxYBAFE8QwfHMqSzceq2806nqi02XYCX2Rg/
saD+rxNaWP5sfqQoFshJWtgtRUcxcrogRcVtHLzU4iVcOxixEqlAndqeTmzlWSOEUoioRFIKdbIr
3GclaMA0qFCFhI05BboQ12UxJ/+4/4+fpPgLRCdvRgR2hVji75wKCSMZUGTmfIvLB9SqirklHBXR
0ltlexTE6QOFo15fqkFBRNdkr9bi5kjw58ahC21c9PYtrblpbIoX3uNRqfJQ3Vp4rB29yzIwrlGy
HpuiRhS4bd5x2eLZp5McCrKLcfgX4l01fDzdMti1hv6SO3NcaKWjmyV/J6w2q33iC3n9B89EKE0+
BXe0p4sjBoLGa3O6W+4VAtc1bY5t1/8n2z5aTXfM380X9xNOTYY3GgjNOyxm3PoY/h19SF1bcu8r
FM+JqMuHZZ9eC1htS6bwlk5x/Viq/9A2zYpKdaZChdEbn+1CnLyxabzLv5cM6gv0ZIheECYTxim/
6ix5dSXzwF1crjlDauVDNGhpDgXUl1T8grI4JVnyJD8iFHEQa72XtjRXgiAEUo4Rvsxt+TLOvS0z
HgicowVeuZV638o0UZ9k8yMs2M1bObh/jvwv4iaz4Ih2yZdTn0+qCFKlDSTuYd0eQMa2vZCdyYU7
x6p6/tdIKjHNTO6kUBQVJxb4NLUoOEMh5o15Y4TNmf2TtIIW51LnZTt/GxJap2IAKViX7Ij8BzNN
b1675dTSHpmn11B8ajvvyRseHELbsCZ+Ej+5Zv1uR9hg4t/AWya8KhFCl2URiSvMu3m8OysGG52K
qJsIIvMMydMHZVL7nqZpEr7ixJkDq+oHMyIUlwaeJr5Th6s/DcUVAJbmCIG1E3xIACmar5cItRcW
xju2i5Q13p3jvGlkIOKmwNAuJqM+Igd2YlekF15LR5X+elri2EtnEf+Zn8f8EkZ2iY8V5HrddHaF
6YUPj/ySuC2xF6K2xmrCFB2LwOO6gnTkcaHqkIOTtqJUMgHWs73+Itar2Y6lt1LGzDoOMpQXe4bl
IMuZV3OQQXZJBChUQRh3UMMfOgIOtw4bCY4V09bqGkHFWUjHWKrHrocP0DPfPA8T0fxmb1cXR1Zc
/oUcFLQOC1h136o/CP649IXvCk1tK/CZ99DwTEXy04V4ErxcY60Sdn+qr8w5dDci/SeHT7CzqPj2
hv4AOyGHJ8D8tL3QwIoQd55pNQfaESIzfufVSd3dbbe9Jf0Qqlblo6LMr4pB+c07Po9S4ObL2Heu
KZTXCgmWuyR2D8uh2eJD9ubDPdYc70WWj5eAV8XxfjPoN1b8drji6Vktxoi58TD8hc2j3gdgFjYl
Km1yF9y/pDDIj2yZYsu+k7gFBv25BlFJjDt92krp+jcl/3ZWQaHhr7rIy7lvmyxjhEN6STxrn0WA
AttTx6uarL6OaC0v9SrPiRImyj1yBberPp2WgDbwUrBS3CWBeazCeT264o8fg1VrwCHsgU4rY1k2
4ZBu9yiDviI8IHiH6VhPVLGrtZspkSYG7EhywBC852R+ZcOskJN0JbQcp/aLCzHdUqYz17FI0SLF
8mzNnKHe++whRX13RJVGmdezLX04VMRUY5+nbKNAsiTwTTmTVY2NWhCDaV1svepIBaBjqEOLahuv
XG/+gbheUof/bgVDddciTL8ZJ45AIcQl9dvT8Iyy/dj7vh6pNJMnzCP0px9km3VB2wWlVIuRosJw
2Rv281kM66BGQlvhLdq2kOHXJJtays50WSlmbWQdoAtfy9BAbGK+rvQOA1yvgNMi9Os2FBKg4v+7
r+rY+R9/KgZyWxcITsr6d+B/Z3QwdlvqcTNdgfVYLT3X273ljgORbR9Nhtcap3DItzR7d/4P/5gt
Ni7dsDEcaYFOonmFg9nsvZ2Y5jlBTcPbAE8qkKlziLuggN4BNu55/Xf00W2vGQJLpP14Qmvi2h/c
HKBdRwFErj+tXHf11YK7ffEs/zRpBvEHuGdOq9YO2LA3cU9NwBzY4u9eal98TzRE98j+Z4dEL9I1
vel+XOetKCLGq/ooAmEk65QGBef+KvEzmuHoDvnwZdVtSiLr3dnJLnX62oAEkklnZIMU/kL3qSzl
4G/yqt9GpKHHPj6kZdIIQPUGb3GNH6ipl+d1sRHF1rzENiYCwahedHrFEtP7gRvz+Z/4rnKkxt0z
ebS0EylRNb695Y2FoW03kHfMnpuav5+rXi8BbKASp0SoD73PEi/d+J+Ho6/Uv4i67YUPYjCQLVEp
IuCXCt5TrkDUCgdePI2QJQfA0CjmLJJ5JwcQM9c4lpau8HZ62CSyj+pgkBPq75fv2CqIQh4ycyw3
EwlR2Sto6wqRzUBhvYqmonOWDcdLV7EN9tJOpMnbF2RX0jcB3+ricKOPSAUZMlvgbsDPd2ZQZuSw
7XPm2TUneGC2v2oF6B4PBHhN8qemHhnMp+cNgz0XaKVM+FM8objAIOp7XAvSgzQPDCSNk8tq298a
1qQbTncE0wwTE0fUc4dpYCY4lIyzCobKVseMfwkwVS2wcXFP5m+eLfm342l+D7YsNt/norvViVnp
kkTZ0i8UQdqmUI0vgTnfnpabLD2SNHisaHJPW4kfrJqo97Yw4C8s6IifNlXoVQEtQEchce6kdHEo
O3rz7jBipegYtbEtPXQ8+iZwv9pix1ECRbTjlN4MspUEdXXOMXjSyOpVwkM+GJyU6XGjMveHe/VS
VErY68Lcgp8eSpuQaWYLkQSpiffkUMBhX/aagW9YT6awlvmxxuH9+XU57aiJvwOlYzZcMZ+8tBHs
xfSrojYLv84++YG7x9Oh63ytGjMyHuh3+ILfGSD1ASaGOSttfST1bQjXjZosEtyf67nBDC+8KMa4
LWoXVw/IRvwmkBPYczqxfu5HN1OZjcjWCVfqqT7k/EXOn9fdB5I7orCepm8mVwfgrNFR/wsKb2EB
d7ramLlJWT3YQxyQ4WWuNIdht5IjXuvPkptoek3P0P39370wZ4FwEMJiU6ra7MXKdKvYntEROL2l
UYeVfpQgyJN07fwUd8tLsLBqawJhfh6IryoEcn/tc1bmwkv/WVg3o9VVnTbFyXRqTUl+2jkzcWFx
hFB0DoUx41Fpj3yMcE6MmLJi9HlSlm7/25oneCC7/6VHbPAIeoztcIZo/c9WJwpWSwitRdMAkema
xoJyvCp+lWudQvxjjMck6hzlsKEUsAqArF1rnOrSgDQQfDevqokfr1fEaLm3YwIZriK1+B/qBx0O
hL2R8MbXe+9PDc5AMdvh08Wa48BSurBwL/joXVzAdxw1xJH+FJBKdbQzTHS+Imavey6VWTP0LWjS
vzsXoIpPXRc22WkEBCBeB/dPzMDIyllmZ7zi83TqO3NlIrYmOQo6tsgI/C0DfrzLa2mhc6nXhLYi
/uiz0tIRlAvdQ5z1xEjW1AYN/IIwfYgSyT1m9An4ujW2bENu48tiK8Q4VU8Cd2pKC42WZUaSXFLL
SqOiIQ8MeAST55N6dPuEbh7w+3kvfRBvYeVyQhwLenEBEvBPyfUDz5boD+8zgSOZLkcNndzVXAmX
YTXvXU9wSJc4YZ7sOg8b5oG7UAEEviOwguyBJAV7DV+9QIbl32n5Dm7zX0r08UjGO4MIDhbahN0t
f/WUQ4wtnxVN+W6d8CuuiL3llcz7sECLsvRh/I6A5csYIw0+NJfh7dHdCH7JWHT0YcvTUy6A/Hn0
DUPqRJmv++WHTPoq6YHFwjWs0CBYY/C3YlDsELhCElIcgk0vkR3vTx85HXF9WvYnfRvaFfgNR88Y
LK1JzoTDlcl3N5TyrDQSVz8HL+H0g0EeSDW+leYHmnN0Pn/eRnPZ6urayDfSHkQaBQ5LoKXS79Vc
gZr6RWj0OlLZ4sA9hSfnxWj+0FzQjPPXm9wa2R1gvqjepzLoob/BrIcbEN50u3YDwbGB2gPORDne
EwZlWsq/nzyflu72weWyjNgQ2hXNagR386I/m0LIWRamYDcrgdc2JY+xRFxdWVqFrk1s9VrG99hK
qduuA/stP2uHByIdQkIDBiPPbue1/svGF6+M4bhgvmTh6f9/Z1CoDhnYcq5WRfzTYRJizTGZh6eX
zEK+k8HhD0VHxwH3pZztVW3A20G6RzhJciU3CsxXaz0qWJ2Qf2VwR/ZWRJjcOY8UUEzEWI7eMvHY
xxqkS9tKZ/qqYyWKomf1+Y01odbK/cdX2M33E7jq/4vnvafKedIymvVxiC0EewPZ7P8GdYFBuOc+
IeIboa3ltMEPYNgiCLPePD6Y/oVNjoIukE7SzbxSPE5UTdAgC+EgbBuHEOTe1dvFii8Nm7Dq6Zq1
YhGN6xXsTENG51mksmgMu3nGyTt4mVPhrY4+FdAq+ddJ/AZbBgKr4Wp+eNampf3pfbS9XDlbRQ3U
+KlaZLdhIJ6i9HNTFVDuyLn+DmRnVo4BKCMuDRsJK70d/sVC10qyDhvRdVs60bA03+xfcKVYRK92
g8+RKjE1f9An+Wxr5bL/Pfomy2o06GajsIRIGEEjQOf4dSp7AZLGK0l4YG+GO98Uez7Y1MxcvM/c
Tan+SgaRWlDh75hRepKRnuRTNM2svA1iHYNUv4ylLzDfp2Uiyy3GPl8FZLoQe9CAy+6Yd3tTIhQH
pcOTjPZu8aTN4eKZ5tobrb9swO0sWCDv89WHlvb4kVjv9kcVC9UDLkMtK8DpyqEuCKxEsaDmsLd8
1lYRvDsZnlTQpUZmvxJ19cEyzp8ClgM8mVgfoObPpFO6IgfFL2/jDTsBudNSuuqj3TAJl31kN+9X
sgB0CxOBkNKLLSIjpol+iTNe1guwAdScflsQb378PiCKf2U0m/lWM9SYnurp9iSeJkQHnq5SDEIh
h09PEx0lJyOA6b25dNY3yuVqI7FP24vFE0LBZese34b+Bjova0pFWliVVymIJzbXAuezFdFsxRey
qEiNT//VA6x8R+fuCgGzoWX26ghKIojcBsR1RWE1Jg69n3yhpMwiiy1VEAs/1+O+xpPcn4Bp7KeI
RhcDBR0kRmaAXnc5KKOyfDQcOBxSgSJvcaV7qwnM4aTOGvHtL/6a0+gUNEyxUKnAOnuQvMpVwohZ
N5IzkS5RIk34cyvItj9Olx+8BJqX19Zlgz15WXZVNQm7ZlJYPFKQH5VQFYHAkeoePxSbnOXVvxEv
AVkSwTwEizNP8fh9WcQz1ce19rsxugHbODXwOjz+SWQGBC4/dnM+6Vu4rIBYT0QPyylEuJiZ7fM5
WYQzB6gOJnriFm1eAOEUW1A5afSJcZprx3wbWBnOE8uD7q+gXRigjm7ssYijzO6giMYb+rFFjad8
EnEXVzYqmAOSAXhf/40uoUjPuSfAUAVVo0BgrYJvQ8eCXT/9hiDWL7sTW6QpJKIpF81gV5Kw0qp8
r/wlktWMUwC8bQhn7RWrH2HpJjlkZnVjpEuIsEnhw8K1SyEZOTb7CWw4/zL0+Cu397fr37LFoaqW
/PDCx9uVtllWabqvd7JRBzgcZyJc5HRI5O6UTzGXO+mn6hyur7NwQfErLpgzjHp31bYlDOWyccGr
bYs42QJ1yWL4VAB/JntgWrnMYvbG+X0DtI8+ZBf7Cyk+l+c2EdcJ1hAUI2bMfJGdl4CRY1HYITeY
+Vk90aLH6h0YUgpZlaZV9HMTgQIZN7JWf7fuF4AiuThHQTohDy7nV2NWWscmiNDnOpA3OL+XCXWy
j0XjeZGzJyEc4hp2vNEOQchbimSriWyghYeiJp33gCDXfr96ptigQ6QcmZICHf4wdt/WxYgRJUkR
2ZuintA25kHwe4ivbM+chxHZFUolBqw8jtVS3g+jlFOFfLDN4dz3SEndfo8xjjcOMXI/GfUjlUyg
esB3Xe/Q7mwY+UsPGIog2uFEimDFdabp+NFQ5mIcYhcxN9t5rR8nOAoeb6bwDyyXqKVPCsRsPF9y
v2oGrRuc3TVDKwDPKjgxo6RO8SaL4TdJumoPQ3LYQi4THEIZW5xk+AxDrjalvwBmQWxK5+82jc9C
ILenDBhDeqwFKl0suTaf0uwwH4NeYSSQ4DSulsgbombIscyjUEmZxNFmM/5yitsMRlgV8D4WcbEo
DHHiUf/ypltDlfBzc2UbpSyHNg4EijultnjvNRRDszsKeqJDN/50oUGLI/BRvep4nHx7q9y9hlNy
AXct93NjIdaNOzHW9MF7zZt9F3dy0Ux7qd0wiiTWo43G+9h4RKrKG5wUcBUBvsPGBzy5b+JWFBOe
H+ZI09gcnADMOjzxWLPc9OX/4ApEzyG7sq2imc5GJHzsUrDMjxUWoxPkBIqnhI2tsUtPqpxYOxj/
ZUrvCXP3D+GtZ71QmdK7oNr752mBR/IwtH6ohWMPc0Cz9YRkkfTeZFQcMu3BkN2l+D6cr1Iq1/26
O/ICi1EARpoZLIQbm85nIjDW/r/G3UOp0EhysTJS4WoyptMF+9VMmXzSvVKuPaeZtdpGnNiEZyqN
GoqLIpwEpXoJSKOXvv/2dOzGGdRIBeW+ueCe438T/CYAC+/Gv+OpUkx2Ypm7y6EIdTYDgB5vUMis
8D0H0K9S0i4FUqAlhrxUJZzr7PJp8zl/ZWvAzv92bMc1jiLuTO2v6D67EmwncQcLTZRUgro4Vu8P
JPpKCUE7P5+WNNaWuo/oNbiBU+v5AgtJBmqB0QCJYgyNd8UxDQu6E4OXDuRL68pqyW/XbDgWlrz6
yjzAPYE9ppToSrsdfkaCDCM7ggNvdtVSO3X/Gt8fRKl1s/uX2G+Bct5+xM9pO9xJ3FdyZ7oBh3D1
BNltYtKn8hznlpeS34IlOG/ZaCeR2m/pJ14CoSYxHHrlxuJDGXlH3BJjxI2KnzJ2jT1uHHA/qvRS
JHMVY33UYzwGPNVst+yGbN5TAXLJQU/BHcKb9CwMUZxJzcRnqtAjZ1V2sJKnkFrE1kfk85TkiMx4
WiNLwv/W68yCyKdFIyODWyQpgjJvCpUROqMFeiD2K4+fBjgvBL2WQaVynzHAozz6CHA8nWrepgG+
k6zCidJPvrf3Q9iRBLRTvnnDXywmNdjzNt0mO87GSIQAY9QSguc659n4zZ8h6mKlknGfQv9BzN0j
wDyWK++9RNpjsk1jYYezVpYXtp0INemGg5gTajuDNOyDYvCd8y9ZAnW6UOYxrv65jSzIsiMv+GaW
wr/i2tQz/D17+k5kjrGaLN54r+0xAfyt7oUM9jEGf9JijpS90HvR0ufBxNp5KyrvR0+Im6jj1pSP
SGthlncyibFPvf2kCVZF+BXdN3YvSPuVSo9Ho1hWvutqWmMU17l8qrkC2s2eHMj5IGyiC7u+NFPn
d6tQhbolBuBBNAo2coajRbZEunf/U8R6Myu/gNbxYXnolMsqJZebmnGNa0DuUWMNOUbq8inf6saA
hSsZgfNMY0bxYWRguYztvJ14oSgu6IOgfNJd5BjA0kv7Uevl9FO280bszDF3uWKEvj6RvgMc/HMN
5PcCQqINmubWOee3vu4DIoa+wN3nKZPBE/4m9eT9hVLsbHgvuOhy1v/2h/UhiybicUmq1s+uekP1
FmrRxx2Y8jp4QxYNh6a5HDv9wLbXMGkdfOTmIAObq4Rxp05tvr9qcZJzIzbw6eSxKfiwILZ3wWvV
J2jhmDkHVm2NM7ngLthUrc8vZ28RdGNrXmSh2eocSPgqy0HYaGrooHYNQ1Gj9c+PoVoG0W37Igiz
gDHFNKngbeO4jzIwRw0beD00Y6vBuPh8Qtu6OzWYgpGU6VYi728bN5uPUNj1HwPPV+0ElqE6kwor
qe4B7d3nGHFM/nz/r+Qa1Z8gQinltWPEd+tviGzuLkxWTTwwbarsxyyGJjD77I8YP0wvKyQNE4NM
AAhfjrvZsU149heTSRqFSnyB+toCM+gYmo91SYYjib42TWYqVyx3N9D+qSsCV4tmkeNyZptnOX4k
ZD9vNqNZvVgqCSxThL+ertdl9hD8GWuM1GcyixfNEbQext2Mk3c/DDj5DcJ3h6tH8KKspjHiAj0F
cDdiKCf9MGin7UV/4Z0Q9UN6aSVNrrbOnC3a1g+Q7mNor0fajiVu1JWveQnEgL9XOgNXBdwNJtUI
rgrH8g99tDJxaw+oPvfAwwNS4h6VJm76QMNRGcFqbFcInJTht0QR6anMHO1mONW+whdCbg4U0OVF
Dl/PSH43JPx7AS9di87sw2e+kBs756kS54mYTN7/IW+DzopcLUMxrjtbUyPeZbs7CZez5XPkfDE1
fIkysIS/efKfnlpWJcqppmOcQ3Cn+dnuYkiqbmxkUK3T4NdTZ45K+JBryLFGnOyxJi3d2mP2bVYR
z49KgiF4pns3qYnQeXwBQodwi3jPDo5K0XQnAY/3g38NwWzafkLP3NJ7ZMKdzFdu8dLu63tQYFPe
Xr2yB+XgGmvIKkTdkq/9im6c7zcoAKiD8sGHK2uf6TaGsgqo42p2Rukc4T5PxCmwv3aa4MhBEZ4s
WvZHdi3upDaDUOuLHA2YPfl8akNMjsJi8FBCe/8F89NiA9jYe8YqA6k9BpixyuLENS+AR9qaeEdr
JKc8a+Zygf4uUFPAz66VWKNEPphzdKR0Lx1fRysKigVsf4IGznryX+bdLo1A/B/ojXsPZ2Pxx+JM
HHA0Fpac656rE6JVvwR3nW/vrDCjtZioq1hUvnRw9v+Vzo3OSCBXqugmVmQZpoP116AzWI9gIigv
f3qXvNOvcpY5LYvkU9sCLknu8N+bP8jN+1QWSdw5WKli0hdGXfsH76qAv0OKOoShmzrwXuOmuHlY
RQVLVM+MbdIVDcE4KuhIGLkWLYUpq9Yc4nZMn2pVjSc0AC78kgvvvS3zjWBJviFqeBpPS0NKAzHz
HyakVQPhdJCO5bPcPCbG2SLNJRY/LLMjAJ8FVSxCqB8BXiD+GuEjAK4gcBsBi3gNCILC2jFc6so1
WybzqdmCRNotcknV8OKiPvSvOcHNE0qbrDPjcPWvZKoKm8qEMxevylT5bzWmgX2jB1iweXeulV3V
TAE9t3VJvPpV22yktLJ7yCsAYaKxgsn3XnYRlAHIXFrGubFZMQeVd0UMiOT4f/yIjgMp8monpzi5
hctCz5PvQ/uU1hfcxc6hs9WJS+kRRfWkXGxFagdzCpCb9zEpfciGO3f/IYiI8N5wQLagdTNAVVeA
aW3SJFXzdOwsc40Vg1p8bvkZtBG5qOpex6HoOmgdy33QYemmsf+fmS0Rkh59aJMWrSYtVtSl3Nu+
gaFsC0uo91NViPgOHX9rb/PgaBcGYkCFLjbNwkW2Z1WgwFO1po0xC01sRinhiFXqKaiSjtXqqTWw
zUAFex5jVosUTGs48jNl9lB4sMMUnS2YhU0eQakTCI1nrRbq378997qndTQYRLWD7pbpxJgGUV3S
C1v7+6s7u0/FTAxw+j8OisSLXjesl2ZeE5dLs3rwM+Rv3b7nyV9sVq9NqWSdBuLWoTbiR5//yvZV
YhLr99OUNgyFzit6rYJLBQNDyj5iGZZG9f9VYjlM2qJvmiYGOnMVH4rBvSoTLTsbaPqB+ZK5We/+
V5XuT/47OWz9V97F80T5wAr1zL5L2zu8RPZApx/S/VP0NoSsl3+Da8gS+/BaRuCULPUk7JfnC6an
PiROQtnOLxnQiiW+eV9tL2cfdhRDm9I/4cBTY0SwG81j37HpJYKDstkg0bhFdLwJTVaJg/SsTiXW
cmy/RX6++G1TLqrPdvKEQf/gSxGDqkxxsQAgswr4LjevnjvLTMuE/X2MQixzpheJESttOrNev2hl
X+smvZ9EHzYQcSzwf6VFK7Whr8b1+IbFKEHYqE34cGsNtHQnQA6AYDmo3FD6ySU8F3AqcKV/QxQ2
/YmRxIDEYHof4UhsSjCtjJI0g8Yskb/mbuFwBwMn62cF3rahcSzXw4cG+aMqzuq1LzaMnh7YNqwm
J2e/zkkqv4u4d8RwVZ5qhGUWblTageI/fn0TP0l6vxBe8WlBBu8SAKgKvZMqrNcYnv8o5pbZ6273
XXx028W63i/ypprmoBTBozGpGYXk5fuPVPMixhpVEQnhepemKzxZFtzWhhpzAj5T2SBRbfV3bn6y
uYNiHkTXOs0jDjW5qLwJsolYRO1Ak27bCBWtpL2qrJKo3VffUHHLgs1dmFpXGkE5JXqXzsNKLN4U
hHjLPORBtXtmjrKeP2j6DPLxYw6v5nESQKeA0r4InKPigpYagUXJv+CN3/+SIdcrP5/P62XuaErw
+TD0hK6pzhLPSV2LLQus6Lx9DG9V69K6y0lhzpJzrHsIiX+Lwu5WO2uxaN1WG1baYWaAJG/fFXXZ
b4l9kW4vlZJdBANWzhDB65plmN1jGqmZhd3133vIWjEvp88CBDTGBNn/5d6RN5tMvMxV0Wy36dZL
WSj29YnjXASMtlMo5Fr1nx/5rGSRUZ1JyFNhalYh0vbitSzErmm6UaP+683a6QmaGLfUfLc4p/4s
6fZhkDv71xcZQHLDTM2a1HxczVY49kSO6RagD8JRDSayw4SdNjH8n6LXV3wtNDxRAI73iTE5TYo8
ALYqCkiPrBX1dTV9QOeJTETqaxOWPoiHPC3fb0jL24fV033gd/EP51lthZTbFNq7L08wqRvHI1Lu
F3vYiIL3PxN9aCY/
`protect end_protected
