-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
GFQ1RnxKlIVX6NwHQrZddPxiddBBecjkax7VVvI2b9FHYPIaoB73XdVdNDJb+0qtG0HAIpdkuKCC
L3HKprWSFlQVnX4x9VJetSFmxIplTRokXA+6V/5sIfO3sLLxMoC96LCWqL4FPZAdFN3faVpPAlRa
acMjA8oGCcw8Vvqm7du8yWGe4xFmKIbhuqG1TnclefHkK2Xw67V/sSDIK4w3ykDwRrBpGEmScZPt
s6kWNP+VjqEMDzGCtgksbuv1At1HDCW7DDTyKYzmhyJlcEobQi+Ng/R99HqPqvJIZslxOd67lSHv
UuPeePJSVQITSqBqIg7hxuBn80cPOMQ2cIaZ2A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23888)
`protect data_block
88HI/8K41HbfZ8Xtg+xEsNzZLOcPTl8TNeUbm1RQwttbwERulh2RVDDaQr4GneOnvW6Jd/Rddgh7
mCImBMVI0ZIOYkGQ1nUJJUJcPaxqLmY94UTz5DuWSJDkkwPTe+96SRMDxYfLzdrBkwNCph6JYN5b
uotnNkk8umICgEN+OSqBVc+8tBI7y5m2U4G4o7NUlXGNsOl1b4FvLd9D8Wxe/kC+d9sRa8FSHERu
ETh4gveaHgJCbJJNgVfNlhoi9AXwOd89Pk2rdFLcITIGmeZDz4ZPkp9hiTPJtSuCoO2ovnWNUbRC
d32p471WBTYL2dwvVW4e7SLBkLt12/izWzOTxZBqLsIFK097V9GqrKEkhSoIjSakwPXW2eBW/fA1
kbrHWaVJNwHlChjj7033CXIlOdW9E4RbZSZKrfgTwqkybr8RfTq5j2qygnLTjGKd+ArsH+F7O7JT
lE715tiXW1R5BXpAq3KEaxuYW3lFt5khaU7WZPYSooB9qeskKSDqz2PkkkoYNzP5df6evKwWggCL
8VzK2BBA9wH+Tu8UO3sU962MAwJTZz1Gio3a2xSq9OinyyW8d6zxNQHT1pwift2kytyNFFAaapnq
ek1g32lnnSdJ1aOsleenEVGSQycYL90ZpV+J/DnaDXJi2+m2ySc8Mv4oA8m3FgOfjZ02umzmhWW5
Nhmy1GMO3uXlaeYOV4NbbXh3+6d/CApJYgDG9r2VBVz/1+26asX5kUF69YoiDEbgFgf/RY3IO0US
Ws/T0xQkgNIVoJx2KfO6KQ0kAbx4bkC2xuuAIlqXLBgEqgS0Fb6X66rnUxDYMyLmtf6GLpjFfeGe
CLH4K1mrNVkkzh+sB+JbdLuiovM3zqXEK2E8lZH8B5nlxNBYyTM4bcEtoYIxzknT5bw6RodM7LsR
Co4+WYTAG7xPHot/NiLfUmrAkoKk8ZAwmG0CFhrhLrFF4WOCxX+UI6/axNn0cDFuh3vJKWkd6NcB
t1zUVFFaA4VDosHyE+95bi2ggYa1rfpfR0PTiPnScRQIjaBgpbRD1W/kP/qyJySMjn9PMdg6SsKE
D7BIy4ig8VHezSj6BVdwenyiaouFAlDALiEbhAiRhn0jfrHEwRAr1dkv0VqDT4DDSKUpAlRTIC4z
G2BSUon+Tb8PdWT7Vpcsd+AsDoOct7LpY+qv9c4VG62yNqExzL9nLRgiNSvrb/mRyQgYqkuvyLrY
mWhP3rLocF5DV/L4nellb/KrMmx5g04Xv7CHuGjtSrzaV6bsGnrZVH/ts9DJGkhpU8ReOCZ8/hyb
03hr2HtHi2WalSJBfkI48DRpAVLCt185sulHKiefdFvs1qr4IohLwdtg9oaoCiVeX6Y8/+tysPET
g33PL2PTYtakYjxb8t+b0sTNNCCuo5I6NoTi42ilJx1m0h9OKObGYvfJ93rrjWDoSdqxKPRTJMCM
wTPMOqX4nOwthpWQGPx/6TtrHoTRUazsJkveiWtP/jrJe/dQ0C4h+D5Q/ZRkEeFg7zXIhKt5ezzK
RLR2jefbZCOuuy6C5ceQYV2SCfKGmpyp5e/43MZs6k3n/6iuvcjUMw8YYHXHcHFQmJTly57UTt9w
VzZU8aFwG34q3Z7djzoAxiGAH2UASAPHHkdWpyhX0eFlrg6P2QLytaYTXrxXCEaf78V/b11dT8Iv
Ez/a2+1k1r4XDM7t3+/00vxP136mK42HCYxr0y8bqXkMFpfZ8BLnsiwX5qsYMvt05qGo2uNSfWX5
n4hUJ/26rqhjUNTBAlUMtTZIbBZGn+gLlKsZg1rAfqjTpYmsStudrS6uk6EzYxZUwlcIzEXmb5C1
vzHVri/jV7KFr5NmhjtqSBLpcG9IcP9jTbPp7khJto2Pf2DjHFZ85yEFbZgxlrKiXeAot2mZhdS2
BE/aZkvLmZeDE00ZicAdI4Fnz+aQfP52GU0YCpFF5UACdOElJC6Jy3c36tJlgEYv0o8zZ57O3lfo
NWomOaECbRoBRqGDwKYET2Lv5DpnSCqS99NIVvgalNBhO3NF9K8RS7n4cunvbhn4MJMhSVv2u+Tc
w9RxTKyhK4rt3NxCoGBw7l2b17yC4gsjqgUm6C4+9Oxks0MZYbeqjVMiinv/rf60Q1Z1uyAdJtRw
ym1+/dGpm6XjKKDXjyLwqDwbc11vMdnajULpQjMxjePuK+WJXxXaaz9YPflp3AkhcGs5qh+37ESf
uVBEuJJu0pczgUffsHNrJ5cTr7PSoDER3fHW1z3SG0hV/nlnzUvVvnXT4XvDozVgty1pMmhZWjUf
iD9autSvGGBonCfYuz5jCeEjSynWnzvy6tO2WqG+KIPmZL5M6c+ZU2mvHaPmNp9p+NW2AQxEToAx
cu1J7VAV9QZ7lQBxtK95/xINK/y5LDtPyQ0tAcRKHAkWceFE4hq1WI1/hTcF4YL45RbheWmgewqE
RCes4lfPPuXE4Zq9OQE+Bj26IykjfInJx/HIV+LXgR/ORwOAEjHAvjVo3BXL4CWyENUedS0olQ+S
F3oqbNwHDU6nxE71H0jGUvOoKKovKA7HHRfCveWIS3LvmSq+oYjEMiwWK5sjXGgzu6Qbrqd8YtF1
JyCb1hj3cSjeTubDS9Br8kAsynkWW91VtQ7UrUBhrlcSS/VY/CUt05nFPteEbruuDdZGX6Hd01bl
cMB0HGEmCdCJtwio9gprCssK6wuh4weALYTmI1fZPLfHYCZMWth+O8Hk1gHpVPsy7z5maUQEK9aT
vNoAIPXvhdm1SRV1fmtd8GNAyO4vOXXG3wxnpGFix7GE5t6fzQ+m0/nwzBejsZka/MRz7jzQt98/
7HFMGKx37f3C/J+08k+98xB9ydsiIKYv6DIyo26eMSORuajfNszjIMSeoC24w3SZFxbRJpZfD6Qh
2LRXgRuU19fVJilPP23318jC5Rz7ZlUeZwobILp+S3X/nBrkkdOJfypGEXybkq7ZIieDRNq6/S8f
FaCYNTgxdN9AcEmLIhUYOL+5fHgET5kxFLUvbC14o5/xtd3FhE9WoNo3rElKGZ27BxtQpPinKTXk
enzqN/6+MURikcYJD5R3tB3kHuu0Gj29pQQcSL/Ea/2GAzYvpI4XRFqiPsQIlB7yCJt/yzO47aye
r15X4zcbOmpN8ftxY0UADFIaLOrH8VD5SWj2Ck7DtIEEux5tb3E64OW/bFHumSgb2s7uE+4GRtK5
959R/3rXFqRyvRbd+3fGQ053mrHa1ZodOkFNVLiBezcHXW7NbSB04ZPmIXdjapZU6Ij3bgL9vQ2X
M+Q9/4hVu7rJ49B5lXvdzJ8NFXNeazCiDTRcU+GiYSDy4ekkSVhlI72l9dPJqkx6MFAr8cjWSkbT
vfvEDpK9prT8bzFZGRHf8veDSWtL5/8vPtuTZqNUyI3/YGsKh4UKE4Ldmj6NbtTmt95NDor7yCrv
tWfBXpCOHE8Mbsy9GGsbAjhsRW6Zodoum+CFk/NqkHJh1DRTMwsrWscxaZoT1SuSN6HVzUFo4QWY
w/qmwDZWHHznXYYfHSixFHyFEn6mSzqnHCuV5qMLirq4O9Dpna1YPNvtZxgzTr8EpT15OI9DeEA4
4ugT8TIQyvxdoyWZ7cGkiwj2opNIY59D2K50+z48KM1sLowkpjQDb5prNRjm2yzE0rvmoSxrXspb
ssCIdT4Esa9kaeZ+KdnSbe6QaH5HhKrq0dGbIAiGyExebUN+bl2UOnZQB59dxMrf1cP+D+gZfqgy
aG5+1K8xO+A96kb2I3l3MAAoaQIA5NI4LBqLq7jF2hXkK1UUAqh/KfYTbqvtwo0dtUG9w+Wtxt/4
mtTnLnm0zpQpccJh2nN2ZXm6luMiDLIE/bsH7mQKGwifLMKtRqJFSWVcgXnQQn7CPLIQ+eHdcA/s
/0GJVlc5enocuwrI8pqoLfnbKB6rsGvPnkJ0k+m6Y8jpCPa3jsHBVkGI8U4YhGhW/bX114IVT+ns
WukTxSvrZypigo2xjhQ2AZfKPu9/7m/PV9MjEZJW+Hc5hJoQlfXu14YfWJs77+AlNTX1OBNzrCQq
UH3CO+hs9/9PORguBSW5gcdyXPmhk9bXOVO2nmA4TmnS/oaWD9bCr+EH4vh8c8nyeZHvMgE6IZgG
NxuJhPlT+M0EU07jt4l3sEAPlBNDLrcPW2HGffUDQYJu9iQJyltDv7RiaxC5PyIA5lfWb5bXet09
aJBvHpoq139mFBZyxmUHu/4ECbpxu9+BM+I/rVjiob0qbElXGn+w7LG9ARtp50O08PzqcfI7OhCW
hUzxf0zt21ebj1kU3lQJPudiS+Z+AzSjLIAQrEtRbFkYc6HhY5rQJBr7XpmKDMaAuzjYTIwJpeU5
Mg52P7Pb3V+5F+jET57T//AvVOJXsHFbqXn3FIxtcuKAk7/aHX5fH3Edp4SnJByCF9jIvCZ2aYqU
IlkchnRSqQbeG8NXPcwKXTaGXV2SkNU7rG/r8s1xsVkLpEU230RjplXBr3ot1iheiSZVzRhOCv9S
rek7aeOVt6yMo3405c3oatSXAw/QvdIZC9VFW9UFJLa7hZe/deJp+9yWZUYpzkLAb4yP2KpuhwUS
s9FwSTmSPMTb0NqHHH5Nnp+VBwBfjY97xabRiafROo3QJLz/0r/vXd66xDZdc6jMCpwWlguiauMo
v3UX72Ewp6DYj102s8bZ2O5YHFjYNr+NWpkmTVtVxEzUBhTGJSgZfx+G0Fws2dXXOddDHVMnGYwz
IrXE7VIHw56u/ouS5rB3R+srdCl2QC/JXZPSqBeLxSukE6AX1YfthdUGSeR6g4EhZ3twCF9rm6z/
JvwmMP0zwfV+8RvBYYLlKD/B0tbxsXaAjJRt6giD6BjhspN4fvyhdE1anIQJa4yBpqseKLllbAEQ
1ZxnmHknZSDoB/Y/ySnCCqdgD7DA9x9hkeG/oEeJmorJF8oVWHsieu68Bi7aSx8VvrcY3rUK4gd5
r9ic8p4XrOWp4EmaTWxL4qrfSHU46wfanuaECYDvY1RWL6VdtSUCgTCrkApuybUzOi1J1BSfUkLV
dOqedaiOvGhNAWMzJjC2ClwydWHGDHGO40u1oZVDy8SYnuwc+1mz+1r9PygQaePCty9L3oeHIgbV
xVsndJbvw0gL8YQN2FsM0o46W+msFzOKhJYnzDwwKUxQvy5327xITpJbyadj18p1EK+sCCSz8mJM
WIjjrv1DbG+I2mRmR8HVMTIzGPQj7P+M+a0KRMt/4JBh2hKbrnqnDUuk4nw/n55FDCxSCq34Bb7t
Gb77b0oewWjeycfOdArTBSXNFSq18x+sJiUE+8EWTiFanZMM/w6QtisQHPaliIDPzXBPxOABzFNW
SWY67wFtYWO12a2GhjBmLnzdj/lhLR70Xkku24NkC5rFjcLnbNvlGT2d2wf2WZDSsu3xSTzmVZRk
zOoWlfbwc3NNseoa1JQR0tTVdsMZegLLmFKQPdgCXhTH58p/IubBPDQCvGYBg7HwwOdYgV7yKufC
C+IjKA/v0YCXEsRdANkw2+rNNNGXPYnI6LweoEg4GzuVtOfBkIRhdSBD8sfmq6vDul4ohuUZq5cH
uK7Ibtp7n6qORUwGrpyXTlDKSA/A9FC0nlaVzEdFDdCOir1q262Z3RDtx9qKvJQ2BY3BE6RNopig
a8WoILJu2bynsVuEvoZ2+kAZ3Kk5MzklBYk6uPMAgZfuusa/vwFj0KavZaZkCueKabA4uBDoRE0h
AQnxptXq93Ereb9mhr16MULGfYSnMnSqerIaDzxNAGJljMeEozSTTGGhyvG0BQ1H9FWXR/pbZ6sX
sMpDNMCQ1iKV1UkpAZE8Y5sA6xbvkvqTBp63c5hVyLN9MkrJW8D8bj0aEw23vyiucczhCyr5Y7Dk
2vY9pi7SZK0BkvipAuqzacx9ULpnDU+yjrOZ7DJg8VsN1Q3B+gzItI+gVhFq9/IXlI2Jj3qerZS9
7m/SrUGsqTfD4LuB/P5vDql1FE79B6bC55Pue3v+FfjCw8iuxiv17ofQa2a9or/g9Pq9ZFcjURs6
N05J2K/STyV/TOcm+D7ef0FU6SEoFfSG87QhHO3KbTBnJ6chVsU4JcXPTiuobkTiNZzn59uB+O47
Qa9Mpmz1uOm585YRlYUIz5fCywJ+jYWGBOPcGdGK6RfLh736G/UNd7+MDg8oeWAtO8Qz0ueKxkdP
ELr5wo0xj077tctvycAKFOcBe57sLU6iEFTeTWon/KgFeeymqAu17uJJj3mXJql7ysWYp629laGH
5U64t6pvooRafOFBKvZbqohTQuz79g2G+CWoZmJoOcIPZj50+81JFWii7Z16UAGS1x9P61o5MT5Q
uauQst2n7j+fhVehWwaLllIqVSxJjsHCmSVL08PFPZ02X9mtg8rDTo8AsLxw9GtHHu4E3sR956+k
a+RZZ6izv5gCToSKZRwMKDMPSVRcYtO9E5cPC8q4zZ6+pX0MM/PKXZ8GpZzvbbpL6TakMJmEQbHQ
6g/T16VrwRvL082I7z89/Gqdk8fKC3osSCPHOJPAfC+x4QO4g0tpzh0g+PQcPt+YThITXGudUWSm
OElwNclQyN8X73v+NXR0m8zgirAo4BHsBsKVsHheTRyYLoG4/tu2P1zwHkE4pKdYNNnP9oECPpG4
Em4Cpv0Zr1RMzQM305BZeD4ynUsy/hRCQDEzEwDWBkadYq9x+kS+ECQYgSdBToEROWmGdUMrAuiK
6TlVfXy1t53/PvL3blU6eEcxqKQT2vj7sHhaftgSSoi/ShoDyDuwl8SHXve7xvAKbs/n/tEAzVqt
aWqV01wIXyxLSs7xWMAN0z17VHKSDTjCdGUKgIJR9LdCmhm4Nd9W7jy4OTAXbGoVSDlR4PfhLsaX
5M/+QkWLCumfIGqnWpVArnP+bvAgaL7QHNAIWeqw1mZWI6Y5ZzAPu8ej0AwyvqfKwYBrUdDfT0Is
pLYY0fX1IHOqnrbcyCrALIMO20RFQnj+SqiUr176DLcnGDCZiMG0DgCIfLB7UQr+mUNIZUREcgVi
uk2nJs3eUUIwN6xkwoJKRARrsk+Fty2LVGe0VUEzTz8B0+cfwzfcyaXUKWyDakPE0+wfe7LP3l1b
nviVTuSDId5dDeXHEYkuVEk3T4j7tkMOds7W9E2yLEaDL6lUtPMFchG++j4sYorrq3CtwbTB0iAP
KrGynHMsBhSixjQPL4ogO/lgl2gTMOUGkBAotxhGcfDKXMRGXa45/pquiioKs/yxsFA/uRYC3wOk
IaLRC6bCj5Zpk9cLAeLh5j4hhmJgEj1cgvDhoCoxdUKb9tuyoIjZqrAd88EUShy44cnmVUj8swhG
MKVyaBef1Ifn2MZl4LEPVqDL6sF9Zwl93ITR0dRnslJMA2E+uYGZqBI8hgg65k8nyvv++1YbHVqh
J5ry4+gPL+ft5pVWKlbhtktndiIpwKfCAsPysGSg4XniOpvRqCpFsTDBgpqQGWENvZRBae/ItNbV
Pl+y0bPdPICwCEQ6o6vKGm8xFRsApvsnmjlohllz3qD5TMnrkd80057g5gZ6Ka2Sf7rkGXnPcAMi
P+cVUXSudtfqBmSFU5+sz/NkCgeRZ4WrGa2KeLFhEPbErMZQfI9WNfq07YUVrjZjbBO3LF8Ebm02
BO+OANgfUzATAWCwNg8k7s5AqgQ5H2cPWTR9zSd0+MsXy9dsxRdOimWYQahHP9k+ffxne/MHjNoL
8f06ofGqomuULMxeOmWiBMOW7+BFNK9EdxFoVkBxtpy6U+W7/ppv1FAM52gzQsM/28ogjUPsxVYQ
ZIo5iuz5BPB0M7NHTO+mgZ5llv/cWFUw7nO0HTqLXGsPgsiRgqXcobDZOeSoZObS7A6YodZLk5XG
ZAtcBdQ4qnSJ3WYKoMM+FABRwlO8UYG6xliYyGjzoN1XFR9dmZIRcRKXyoWkKW57arlZeXv5Ybe6
SeiLGZmpnjKTwZ45XVn7nybVMUp3knGrMn1NSPaIAsb2Eo2kHFuSG3qIbzbnIW6r+4ABuabrbger
COZnBy6QlVOgkgvoI3pxph8LcezzIwfnJh09FdDDkmoNUMw66IM6BuTkLQmqgsCaWqPXtH0vRx9p
pLgdovu9qBCEXwZ7Rv/+1GNoU6nza3LvdYnPI7IAnB+z2TLuilpup+r9p/KXjdP1F07zPZD14oqs
paxgnGLg7YdZeZjJUjtlKvz4rxChoieC4uTfP54zA6z7KS+Vt2xnxivFo4qZVFDLjHGfq8F+x0yg
+DoBB/uSXzaPr/5n9mI3hmsAr221h/4frztzvua5pLD8mctrjEtvqQW1nT/IjKzpuysFMm3ey/hL
csEWSQhhWtIzGDjkuJ7zhlx42qTlamrk4a2/OUG03Gh2X9u/N2SSZi5y7ZoF3/WH/F84yZJGZgeo
TV50HES5n3HsOcuJEmJdsrjNvmJiVn2KTkoy8hj4oqwUbyUqnIgSai2zdiNab4mMqPr4dhM0RRAu
Ht7/UgQutTakhbfcpgsfaEax7qIbukcCCNiKzPkMEqjTpJQLclohM/7wByuuMB45tP+zb3MDBD2O
FH/ujMe4aUtFDd7N6q2wBs6fquFXEEm0joBK6LuZXXgpzZc72vkROx/BqEydZZbidxXEWqdsHdUX
CXqRdecgOWeMWrModdFJjr0CcG2pP2iOKUuaTyOm9p8mKzGVOdZGEEIZZH0q2STwLYTSfMAnEHft
OsacrtVOhoB02R/1b9i372pVoB7Xm9dmawZqA7vj6YfuQ4CaBwfweyBNKctQBuVwU9Xskhgexo9E
mGYWt7OrPBOrcYe2I/6CHYSDBg0ZOAZ/A162yUFBUAylxoVX4z6xy/b15BbRxRVN2YjubyJEH7wk
ZzonHHveecubaLGJZhh6T5w8Mi23u3i+DU6qsPXLA4wIbJB+fcOYYo1D8ZyN5NCc5Y3FJQN0duu7
EOSvezBcq9dpZpnAj5roIs6lZ3pDGY7hHClV5p1f0rWdBK22rekVxlFDK9O7icpGmDiOGBnDhb2b
ocQaC7+AXWNdhyYvPXF5pv0G2CC5C86CX9sjFjJ6fs1Q4jH5O/x5bdDxPgouCBppcSO/Tuelo2jP
jzxUtV2mWQt4dqFN61frNIewm7NSP/4T+iBLovvjego6zVtORPtTpDyo+8xFwSPdwCOCeH+XZbbt
qmm/81JizqoJAFGvShENAujZQkKqCdpGarJ/de6Hu914oN7k1yh8Adfl7aTpj27CG83rguQhV55U
7ZWtf8SEg5jxAMlwgFE2goPIdqudVPVsRW31L5JMBWW5cEvZwpc4R6xrBv3xqYHERIPZ55qSuL8M
xT7QBrCr/OlAdI6JBWo8B4h6Tg1kxNK+OkkRsHplidASUnI4vXBoCi3VBtkeCzO25BDe8FompHfG
Nnd7lUvEqJahEEkZnXPFXKMyS36xWdhZBXF3bmtafZBk8b9QWLfFDMzU5q8uwDu8a0FuT94UFCvX
NMpcRNJend38EAaDgGYR7r+zPNp+M3e8DecQPcGHXtMu50L3bzvNP86rcr8sSmE0Io0/8H9oGli/
G3ko1YjqhLG+G3WbPZwR8LC66/37jlyCAsMTaQqxo1krdQZntChxrqV6bfXTAnP+5SPilGjFtm7i
G+IvLP7PHAX8BzhSrZ45hKvDn70O0OuiEucrFfjlsdTlQnQzSofwU62JqpOlvU7CSQktcDc6ihIs
0utq10fha9Q3ocYck5NzQlrgO4CTHHhp9tCNLZYF2hPRrb3Iu+lPc16drBcgXl08EkT9lmPjde0o
SzypnFVT1Ta8FbIDWiaCJW7BqgNdyi1xzynpY9CtYhATR058NCjjVuNqgi3fZrnzbOn+PR6gD/zS
1LM4L985DAWKxguubD2jKRQsTDEqIEmv7nKoCbood1i1Eo6zqcPHBToKU/a7HH2mOOTj6rYByuUQ
GoQ089gzm2L8fM/G0QJOFeLLFymuMG90oFYg4VEup8HczalrDMkjvrsTiioMN+pAe2PN2Y14vj7s
QtrE/1iUu1gJXtdVTmn7UUQGPBVBxdxOW1fq3+fRVGGuXbCLS8L/84UGcgPg8mCnLkGl2/NPQQk5
lCnHu6fqF2vYqSdfiv2iJhfGxIDYtTSzAmqKonRtbgBspfncqV47zX1/3Wg6PnaMsP/OyMsaWnAB
TAWWnVqDACTDZWl5qN2xB3iTi8bWcZBamh1WRXVkdnWaH9YG5pu8bJ0zCbtWKqGO5syHrHP353iv
+kKh75phnnz0wDcefJjpz/K6tc6fmTtsLUQbWwfKKx5Ra2/Q2ncLyExYo+7kbAAGjsDjteMFSfiW
5xxp924sK+5PrRrsXCe+GngabPFDl1EW4XGoZRPjCTOIUjHzTgLv0Ry/MSE3Xq/rQcRauoLv+isN
y0eu/sG+ihVQiF3in3aBRtf/voI1W+xjMjmiipsiuooACeH9qyGZ0eG9Jqd4if1u6fFTxU8kWLk4
PIeZxcyfbpJvJ9b1JdYMCcdr0AIaaTyYxpsSj9XOzr/8NN9nZrOf9lcXeTR9mCxD6GzilRz/nOWa
4ormc1vaD3BoK0npYf8ritlQwB/GnBcXDxXq6qS4viA7NMc++zPowHXyyo0aZWSDfwDw8+1E/Jgu
3TUlC+umGJ9jImnoTHAZ0Jf2jUzYj9R0upAjyJyVkUcyErasdSrTTmaTRnKnwtM4ba28ghcJceM5
XkSG6ti9hRr/kw3ilT3DnRe1heTFtyaBj1u+lMEPdcvFFarfGLZP65xgfuV8H9HZ5hTIemiBC6Jm
8fYa+eI8+PWmAkMn8wUUNgyeCi+hChcVJNujeSTeAoGthDZPlXIOGNBgqrcIH7rEHUgXUoxQVv7p
MdX+eDaZ8a/tQdCMerNfrrrdPE0eYY61cZRD6R+S0ZPpn9lYQRK8cK5FNhPUhZutBvyAJfSJzlv1
ZY8MHYtXFGzNpsVcIgYBD3cFhjbhpZPmsp7zix4RQ27TYLV5ni8L7GVbgYr78w89dr0ZknMYpz3V
YcgILwBws0TQsucYGqKdMCwMhKj3S+tw+nHmgXM5Q4FD4g/EnRiyF9ehkIlggZ+7/hl5oGUoEiP9
hQIuxoG8GOYPtKheRXMZJzJ9+5/oDuXWzG5nKeyuxUTkywZXAo9hPRBfvx/c7sYrJgzofbK9cqF2
vuFVEjbj1TX76Go4+UXC6pRUl1l/4YUSE2JT1yg1vWH2qnXxpYOuRkRsi9ZIxljpUF1Rer9sB2ze
U4dsbDcytnyySjHMSnBosdnJhKJJI7Zm6rOdKCcX5+DNX/DhZereFHQVYP25gyEjEg8rRNooA63x
vsudFSLdNcucIH31VbIhxNke4Ch0KCqltw5W+GVlFGu8sk/5N0OaRme5zj8/AFYUb5BKGfVBfmW6
khScBeFolxoimK0CrmqYaxo6X22wnsYA8n7X+uBbQUlaYhqqvorQOwgV2x74WlKXZxnuuY3UEZcb
WjFJwN8MqXRwUifKzeG8V5XmRS3APblBS7SAhc28dpf6pFXVWB8yQSMHSKJKv4pjsHQ99MQMAijN
crSuMiMHCYE41LdWiVxi7NFLpSiuXCLTkvaEr3jYsKys89p6bXaxgKoNohYAMQ6RiFdbkihg1Tku
iSBI6AmYT7c/bt4LyYR+/3RccvTYB1KkUWPRggCRMqD6NB6rFbMVtbH/QMP4NHPUqz/Gs8Imm/ua
yhFIpisGQs/W8e5vBFB/zI8X3NPDHKhvQIFNtFugTRSraztO8y7ONgPRp58palJOncCqibik9vOT
qHVHo8vaTq9OPYFRuq3m2eFxuEke7CSZsOgUJu7q5NbYmjOMSYKmu1qVHcqOy2LZ3DKA6nBhyK43
/+nH3uI+UMV1eSvpZBcjVuuLQ29sokBy1B+fpEiafdWHMayXZYTPvyqid9ZjpuQfkB0J7tzSENYx
a48houx1vWADEpf+MtABu8kQg0kvkCkEEDkV0pk6mB7mWeKxwQ7Ea1gvyGU2zT2q+UM4Rli6O/Vw
ReeWVvseMlyUKFlgDLNMESwBqZQP8X74yq9lGg26MQOjtEVn5osmNWz1mV2O37G7BxGwTRFg91ZE
7AcHCAinL3fULWWRfMEu616tMJzH788VDXks6yhKSqqXx5XhhVAmTV1A79lYcDU6rLMRLNsVweWT
12AruckVqbLtyZbGQvc4FdlgCFS/qZfeGNJgs22CjQZ2W5RD/wsrEUeI8QVxfk9j30srmNNgg0A8
xY3Z2oCeG/4XxfZ+Vx0+ZwWvtK227KiX98AsybelZXsbp4usYsA+vXr+u30makN1eo/RSxbbG8gg
GljxuTgjboS08EOHbaS/n5dHJdL1WXZweszBO0np+JX7ykgspP7KsDWTitzIzRuj1JFDrUqp4FZX
bAGYBEPbk4bLeO+AHoHSIPbKQOhWRPGcmdnnndnczp5xLN0uKBuEf5uNIoxV89ZrHxDI/ukCY7N/
0fc5ji65HWayDw/BJsUL1HxNfy2wwxFcg3q22EY8BW3sTGT3EojnZfaW9pBlAk2jrWb5m1fKgEMQ
4YvzszIvhyVkbNt7ihz/A0hEW899ZfAFmPDekYPwaYW3n/NlnZcSSLqJzIHU48C/L/Kyvf40OE/k
CXGJQPWodvORhgOJeEE9KxTX5lSUOKZqS+GAHlz/N7x1EPUot5qSJJK/PouaT/zo32OuRWJOP3X0
8ZW6jrrX3TAuoI6j1w5/svEX5B+tC3W+FJ+4SKgZ9DzfMIvF0o9FxB4tvoqtajD1D00/WdCQo33A
tnY3ms3XmiqUMN1Y3Xh5Zx51EyOndq9/KVl6M9DzfgisLvmgLUumG5K5Y+HRNBV1xOQrd7Ex9noB
01lKlVvwru2fi3MT2sNVzx7E5NPZvoL3Q8KN6aJ6WPg/NYmyJ1MALrx89uUzEPnJg0GTZvqxjuNO
LfQBOKCPRSo8Er3dgVkIZ/xWFv7pNJoKMmpLlrs+BJvuarre30XFfWnniw8OSYGoD+he+e4iC8iT
gEixDKN76IG9AAcmYlPpflYTZXBQtwZiua/sBwPbV3JrDzxG3AbQotNnlatK/xSwqwfD7FQbAKUp
vlBwHCzQuBRJEmLZpr+r7CrUWXgfuKySygVRqVvZutUEIVNJpUhgfXjobpKjpDwaP4OK+NzS2m0l
YXiBvpK1YF+7F0dFMer2oZH5vx4oeX6/sAOZOAjnnqTB7C5MfTgLG/GuN055dFYo7jmempBNFtMM
kXnu2vYcdqPL+xv2LUttRMAtvpIBVI4SaPaBPr24HPjkTj3nqJz35367+pZwb+yub33q3wF/ttXZ
XWIMuHxZiLIwg02/6y06c771N/+hQy4Qq3Ia2aLCKTD3tyYjaSWYTabh6I+nTX0tgUqyerukRIii
u5IP0XNk7I6KbmT1+2IYUMDTBwB1EDa0flAvJvpNk7RxXvPwToIuckb7J71Ba3bGyMsIhUemTcgB
oXmlleoiOZ4gNksUVbVzWjLxyRV+Xe+ucKetzcrxDdvgAHQlPFzUziyJd1Mm2JypC1X7urYDtkrn
sIBCtzQj2rWvnWd/EnXlzrF2eWgre1eJER3zy5Y7X3kKI8YhkhL4TRqVWOtQNzTOypuwh8WWgcp7
atcWM9QviSmMoGRN/HUNl1iS5rzy1twu0PLr86S61b9nbv/taLKS0PkzF9VvPxBPB9cDaHKqR4cf
v0krsb7rTTrUgovrZYa1Q8Vp7HZOnx+7ldZDa5RmWeRF1YkvNuhZvRuvdCpxZKebztIm/M8tn0vf
3tD8MxebyIPzYDjrUCamfG3tKgg62peh6wkRcxv2dDFVAIhTMX8AwJSERqUhtsoFEUJroh93qsAp
BCr3hbBIGKKxS+qXgKi2SWtwt7VOq3Z63yB5Jo+fVh4iBlwOsvPic9wsPLqLt/6W2Byxyj5Y8kWo
EBQrjZTH+MxLFETVj7XBBqMU4HXudSvGPCpv9AqOyU5qFwQ53N2QLjkxzDWrqCVj5Gqel7HlDm5J
wATPvYINGVi3WjolbttStuINXkYFBpLNRCkWe4+QLxqZkHf7JGcGpO9ckVSUtv63hKSSCd+Hpme0
F/9Yp36guLw/iZLJ8aWvhQr0IUbA4VVOnOYMLyRKWMFPFc+eWYhrqtWX4fTNtyolNGsbZ3CNfccP
0ABj8RZOKmMGwdj2LE0arql+v7DfyNiein0xXRQt43tK7jDrWD8t/QjrrMqlKdtmFMKha5RzK4Zu
a/UrOd6W+NvpWk67FFNCXSisinR2veQFCeVgHP9hFDN80X6hzOXqOm0vXk8cqVnEGGzKE+3dnMrq
UaKk+QSmY7KcMCRaQa3HcB6HZAyNjU99MvYyEZxO3cSKmSSIq6txSTH/gbv+iM3fN6Nk7NIMjEWc
C4IoMLYXL7NcJII9yB3weAhFedHUmM4lfXY9J/gw3knMQgpn+pGYxDzJQA1NjYSKu11MDVeM7dWY
KYSEn0qy/rouMxR0/iWoyagTOB8wx79DYnHOSpCSW+wx6JqzN+6eQ6ArUNjxFXT6CCxhw/+QKI5U
Rp77JOATCQ7zGdVF8vx3XlnwxXuoICdlDDjEBX2IROtnpxrxWYNY8JFjpwO7/1LJzp66+XPMVab3
P9Zth+wr1LMGNImv/cawwQ74Wuv6RCNdGtVFu4XE9INq4cbDKAizWYJhC+QlN79QZVkxFKEgcwH0
qrpFfOozpt4Di6NPOra6fqBWFuhzU4qfAR6lpFiwxRmi9kpY5bUJFhgUnxU83hZwezkMP80LwHeC
AftgvN/cDDzluZ3VqaNpt2cRiHIDG6GU9O0gdCIVfBjc+RcMaxP7Jezv/03DWZwKzuzv5/ZsI9xA
q49J/sEbgClIT2oBpVGV6DJWS1oikXOyGyG+JLga01dEcUqdIt77YFw6D1QRSy/Oj1Cl2uGzKROY
Q7NuHTP7NS4tsIo8B7AzLoM5duOc1wHUfLc9+AJDvpA8VeoUGuKxKxPNER61NAnWgyWxDItpIzIq
20R9Q269nNKbsi6UYtaAcPe65WWMGVoeaiddUSr9dM8NCBMIRDtr/02gz/5y/Y1M50cUyLfaOGem
5pBJnxv0WwMjyH/cs89aIYyNb2EhDBPqjpIqNbCz4Cn4lNO3mKbLKbj/0MgiHD44qXzp67kUciCF
VjvjhPsHsZ77QN+/FaOMvmzyKQ5Ouvwwxkjpuei62xaGRk913T0KV4bhxp7CRO42t+5PhBuCH6TK
38qJxpsBJAI0GiVoccpJQ5AsSyYI0PPcHLHkVGGG+2y1qnCB3+4G0+e2Ia7Rf8Xr/fSJOEJEcPOV
U9fIAqrv6XSC6N+4jjBhsQhpPEX4oDl2QtV3iQSZSirpER0sWwB7XfINUhx29dUtW1dDNXOGCqwp
G7ugbAKLhkMmtEuL/qGIw+zP+v36AhR9yhvQmA2tOGgNWNGYTy6GftSePbVp4w2WFdKq2Y6u28s0
j/x0eVfIm1Mz+9ZKcnvTNPJsPyguDJ7AUdWZYrSdirQsP5C2NiMRgq5N1yKY0Oq+srpqQ0UxdtzB
VJxNd1o6b8Jpmp1ceyovf59UfGu6VRsW/z22j+WFUvqe9qjF+QsBMSKpWwTNG0UV36Yh3MC9aMC8
RX+sCIJAmI5wgLDh3gvrCl5ZrNXJ/z3f5ce8BNdY1BqrK674wUNwfhhgeuwRgt9b8LYmMP+0Ieqy
+lDICRGbIAPgDQNBbTfST2vSzNTqdPtfenzskpxIvBOp/X7FcU4872YsT839l2tQDhhOs58ZDpnC
6I5l0C7EGChBu3UGf9wwx2DloNzfiPjXUCKWDb6EEIn0pGtcZGvoSxUPNWXhN72DL/f3COu7TV8U
7H4902xj7Bmtlq/358qx2mYeKivauaASsEAW8xV5jIHt9BVUNpWBIjKK67A9oPDqaLL9z1IaOMQH
UyRNRt3MXigF+eWlG8HEg6flH13OgDL0FwO8/ChbABPzEHXvZ/zjS5OPU6VELay2yxSYzaPKXY1b
rNr15vtbuJUDbmz4xyTcXsgq2bqNvNZUpbviTa4U0UQ0p000OKeg8RhQwTRu+9tY75e6dpMxCh5w
osZUFdk0lMxXt47fgYfgCDDdz4yz8qI/ohO3i4jKWbyKOW4/RtH/2s1dWbwmUD9qy6gj6c11+fYf
VkAoAcxTGhusmWayD+CUXQEHGRPA3Ch21HGSn8XYXbs7iAIFOvk4B/lnI/oxNotX6KFMwAaSOw2M
jSe8yIZa7p8kAVZrhsE5O6H8KmAO+dnZG4pf9LeD3cM6d41JafVdvdqaJRWpRMy8VWz9LKNxxXyj
LHl/Ckd3CPq5HdYwYh9oFkzjz+5vUegCfhefl545Tvz8W/PME8e1u/rzU7gQIZTDxkFCXo38s2Om
M9R39TzLSDQhPWSE09VToSMpgSr5JXbN6O0d0OXIK/xsj1e6IwjUeMbgoVn2a1ZFoYrQK+yLO015
GlNoKjF1Xlfy2xGbOyf402oh5MERf+kWI2GJmDuJ3vK8152lAV9SdwxNPQKiMLquIptK51HwWLXA
9R7yEXJO9MY9ZkbcnXjm5ilCIKcXMQ4p4L2EVBA1TmptlWc1+SLFT/S6GHp3SSLvl+fgJNaYk6Vp
pamdz6VC03nVVBJu5sQIIlmPRTUVZJoBB+3BvS4HxRdEnIVPZq6xcKu/ouomu1SAJmx/JdVWW/vM
R3J/jBwSHE5Cp9i92EnGAvOQ57YW6s2FRuGLKygZmbu7tJAIGABTm6UM6UkUIFdZzAxyUTzXz1Xp
3ain0sTdOgMPduTdRVx1Svmssspzb1q2FGU6/aZD6fslV1qeE4wXJU8L/ZwPyFzzLbFQyplx4B2T
4mJecZ8FXm++any23zmwmZQNdZG5X6ZffiqHM75bTp0F7QEmL2QPC4zHBEYONiF11eFj2oCdxOz5
8wheFTQpH8Jdeh/e9almzDm4oIwJjxRe+4F12ym2ErwK0uZ11Joib5uE+D0kco2szbG5/Sm3gZTo
bl1vEp8sKzAAF2TkUH3KhGTNF4C6zFP/jzv1VD+2Hg9+1j22m1nL2D/kCuDhfPRqk6VXyrQyGN1u
CyS/0EENWOXvLhUmgfmgJ3W5TeBQ8A4Cd4cHup9Z4ScmchtoL2f/GAYwMQ9gq0ekOwU3JXksjKCe
CS+IQa+8BUfCoESpJEKBmCTRZCSihvpUK9dCEMW1gZxxycJGsYY6d4vLq0yHq2kypbpieE9F4hOp
E5KhdpKlsptomobrXix5fGke5aainGlqk/YbPeyAq0THlGzekU1v6loc7+yYncjFERiqVOUDm8uA
TUh41VCSgx1mIEXycWkGZ17dplnqgFUfCg0oyWQ0PdW4dgV+ziJB2rjoJqLwYmvVa3Rj55IYCmnQ
whFHdFjTyEKF0NHyOaulklOLq/hS01A2660LkOm/8s5KWrWIDmw336lq9+8kO9EOHIbTHB5uDXBQ
1Krbg/RE4JVKcYfFZUskJjfHfyPkGecMh9qyNirZX4R10w2lPgYdyF9TmMwIo2qThM+iAukrIWHX
7F5nLFzXV5qgUbSd778Mcp5BqrowuunW64o70eD3bdjYNX1S1aA04J5IIXXBtoQ5CWCNirKf0gJx
YgiVTgz8KgmAHZCPM1p9tj/1vxYIFZeoPxuUP2senz43rnMOnICaA3uyLTZWNcCNaxNJqEO4NKW+
X1sreyXGsfCFtIsEHHbezPmy8rIsH/i0iQKiUxKroHUI0yLO7sx7yElkWok9eWRW/HQ2NB5XgoJW
UxkuIb+ukHvAwWkstQqhOFvHTgxFzl6MESOuGjm6e4NOI9qYkSBpmz+dGQlzjnu6VGxdsfluPvhc
dfaamDFX3jY7R3CKhey0SvFEqSrw8kZ2dEAFeWGQ2oZ2MugBTyMC5VKJiGL1cVgNUDkJyZbkEvqG
xMAm+qD0dajnJOoedWpm/mrPBfUtT1ZbU9SxUrG6Hag3J8gutgsg5tVFcOk50l+3xDR1/RNypRxV
L3CroYAKd5IxxcoWeTlG/dQZ8Wwx8NvV6Ok6zK5cJxCaq/L0VOfA7m6y3uL5Rzh7iws0ZCYzJzaq
dHijtLIRaFDZP6pdqQu8z4z8A3wDoIZ/GWNSYRiPUhkkp9RykycLAtytDtDLF4BWOzqmEghGNWOj
5/RqPVkCbkV1q1FOxNs8HGr/aQdzZz+K3bfCA5v/yoaS/jovWqFxNKzphV6RYwqK8iJEMgAtv6zM
Da0ijm1QPS8XNsbJBaz/29rokgt87T4IOvgFDmksWRUa4wvrn6cKxJ3THXhCvA7ndljKPbYH2fHU
l38BvvodoqYPwYUEdx8u/PTwZpRwbyBc1IVHH0C9PMbzx4Q/zLVziJ6GBTs4GNG84poJ11aWZUfr
Jb7ZokvmQ21P14LNwd5CNXelu8875HkJsCvaljFrUBsCEjDYVozDpVStgermzLm2n2E7aGdrEikZ
yLYToFVSAi6RrNF9gQ0Ul51MV3DYbppTLaInxGUwsapZ64tmEm95Kch8y2um6Qz1wROi7YHgQq9M
nQwTzVzY3gQOL6Dbz9dPhun9gIK8OEkFWZcmlCr4kAWXhxf1V6TfqmN6qrEYL0kxjKjeACulH0BO
YOhK4FZKJEqPZCwruld+hS2PyW6arECiy9X0HY8n+MA52MB640QxQxjLv8hJG0fPRso+7N2Gud+5
HciehKET+5RfZxC1P2fXQzfbevjYJ5bpg8CLHeG0AANRkb9Te0cvUoAv+mqu6J65AhyDxYBtKHcZ
uHbthVYIEv4jGu/IwDLM/HgBuOsHixvdGDwJ1doGzM04cr6uOKhc9qB24bv7glxk3k7DCMxrIQUO
p/qCg4Uaf6ZCq8mNz65CIqZKw2KDCUeRfo9tk9nLX4Dst5pRYsp3MrjUXVy2DrDcwFeKFCjU0d5a
TbOV3sEq7XCLHeWgy8W0BZRpBea+cMLs2T22DwyPdTKIZpAJ1jYlNYx6srmlMQqbWPkSJxpurBXC
7NDmZsGLgR3JJTI/Xnl4IcI1GB+E9l1URW/62IzpeCVfXaHT+aQb3xFiRDtDAjUL3DdENmXFCiaN
0iziiSeB0rCPCCXxubfZCHPVWGVEHCyKVZvhwKnXRFsYgfKxzkby7oKiUGNBG0Ky/dDFMVvqCONb
oPm0/wCvqFCkLutntMp4j4N4RdDuk1wTJboINb+GjpL9V01ZirWiAKsRGM8ACcaxLKpZXZizpmHc
qt9vr68wV9J7pni/3lT12lCPjw+3oYsr2RXN5oNZyFTwBXbpyO77GNy9vJl7d8kEANO2RWcrCXA9
yxd5nLE2btFHcn4xrNFfwAuknYtNrQYQqj9z55lSxl590oYIe3M+wVPkexm0gV4LvW1BDTyTiHQE
rfDN/nM2yiigshznQk1zZDvxc40q771tH5D+uQuA6MDsfvMDU8wdyepwmQfq/Qb+xIJU5TDzTveV
KiUHQVPF33AlFx+6e/RUfewVz5sVNHtHnw+B+0AHplNeAZpggPOr2mxIHRHPseBrvPjY7G4URZ4U
zurZuPxUopcsonA0Cts2gN4eKCyaDKDiJ536WHfEFVyGqRvykozvy5AU5t9/52AVfPrwhaKX8RUV
lISMcy9Sm90N66TvPMfCVOIyDmxbqluBAac5LPLHXDCC6RbWFCU0XrijGY6m36518t6QS39wxuKC
LX/hLOnq9EisIPtENrcZA5v/HWTPnVLQ/SbIxxInXv5FNDKL2ZXp/njIYey9ux6qfMJu29pfwgA1
E0Y/ih5bOxTgF/7h8Ux1lKF84+CatqMa9/t06QsYl9UU2Xtt95y2oAWNidT9h2Qt381D6zBBnoJZ
LxXVEdjXkZEqZDvuh1E5HW1gLPiq2073eNUHv+wiH8IID5eH07TqVuDjIke29pbPD9lWLeXJcVDG
x2NUz+a/YV71v86+hN7sgqXIZqVGQqCMA9MTIkdamhw4ulb/N80hk7yabJrixhFvqgu+aPfHxJnV
IAeQvawRXvTEQp/07oMi8smfHZe9O+ATAhm/PdSWgRhQa+yluHi51k0OGTJ4W24z1MFyNgqK09xq
dCrLg/NAsqpBoH0xJfilGzDxC99iuTBv0k0OwrceHflrAidcTA3K0rjBNhWWdOQP9/D9WCmNiat/
4SKrDLG0oyqnxmRQmxGuBdFffSr5foWTKrzm5MmdntcBP1OVJvF17WZaw5zImCKylV9tobMNfED+
+W/i6LB57veZX/6bt0E9s7o8F/TDsyeFNhUzNYtqgipIjYrUPaGzobRMHVT853DXP1EKIxhGfLLN
5NgGrl1eijmY4B0NFh6rsZqkBcPzsi+FGt2HRGtGDQZlriBdDQyj9g+vWxh0PeYadz01vVKs//md
rr2z4oxsKkkkPCW3h3zTFdWaPreVcs2T46DJcz+/RScwo5f3mEV9oEjcmjguwUz/nGcOjzFnPtjs
8z8qN3aIqw8CTVKYNagcgSBPlYaiZboV3t6ru138pSfwiqsog5e7olYxtV4dnM6pnBo4c7SNbFag
DdZNE+zoyac5O5MEWtQDQUj51nM4vXTagLkhc3ZNG2Ocp185Ef/NzBrcj7FI00PIQOXL7Dhg420M
bCg++7lSOZXKdvqp8yt8wLCAbial/rO1GilVxFK7YOwQMW08in2jYgrPBjiYihYeDGa1sAh/9BPl
3memX9nXxv5nkeAaY3G2qbKXp5HYZRfWj9DM5OTRV6p9C91kAp7RvzorLlTnA1Qw0fB0T5At0Mp2
5KJLGztEbzlupAsAPt6RjUsw5YmL/ClnsJhRScICfJkqeTxrcCSGlb1TFbl0PX54Kwt37Ap64u0i
4aCCJ7WI0r2O53IzcH0PSwe29Pc4FU0OFjurF4xjVtfwoCDZnZceTic6LgyZyRfOTahqc51toiBd
BuJ6T2l9QgThs/Mj67jh+Jv3EvBhzNuVswf1P90IEqK0RpYUm4oUAmeN1L3GJxpNCwlhsTi8JKV2
TSKEJ6D1T4/7xR035s59W/x0BS67ketkSnQy2q1+ikFgupso25m9P5jZlFtwEUInZtsCfO45zvYc
8xBdGP5jWjlNF8Gi3/2eYGp+ZVqel5yvnRYBxHTyCvgpfmJPlOEkn6iJRmWmM1+fJmv4tEn9hyap
0XX8HDJuBpwo0iJwmT75oYfPerV7OUhYP6rN5WzPCcrFg67iTxQ3660W1tmqdJGgLxSWDGYwWRbX
tIBH6NCDdvkDPgOapD2fFarVHl4LGdorByNdt7/oOWr7YD1/lCs4wRK/DJKvu/MsjVaCp9NtAX6N
A6LGVCTmVVq6tVAE+boD3eEZKS1YEFI7sPauFgPmrEq1SJTdRvrj/qcOQ4iqNmnYP5KYDZOSciDt
SeQfaSU9pvhCFG8VEBGBtC6ew/ZMbb7GD+/WAE6nrTMQWvqTb/cgwZW+n1NUKQ7FdxNSzg9QE4h3
MxJEIxPa4fI351qs36rTG1z62wh/v+TBopW2B5vEna28wAiDTeAE3/NVPD1qiTcsMSA4uG41DccS
JMuE+4ELwQRM2KKtyWbBc+8FPR4JHBXsMeOJZR4oM1F4Vw12PIZN8cBo8HnWUbhTqhH4WZaYJaRG
WEIS8y2eGn3gAVMOfZhisYoBDxlWCpLixQNCNV8KDgJZ5HTWXPnhjDriLIn6kGdKZ/52MIwy4jJ/
swgZjsF/VJ5SJFtng1bf3CqQPZJC2+GQEysglGJzsnphvWrWobkNJ3J12Go63dKb1yT9qg4SImjg
6GuyP+vof6KnL0j0A9wqsOO/ICYyFotJ/aMu2S/Lo+Mc41xp62kTKHX+/7BFYi5AwGlAByUvG4nq
kPGjXhnWg8ac6XlEdcMIcaeW+Z/jEHwnDFIYVrTeFiTUSH89ILHJvDIHnn7CbTWLH4QDFFZav22a
gpCxVh5mhFW1RuP/7NHqS76hzz8tjt4g/Um3QMqoF40cyfKZ53OwFfWZVS52+ONqJrpurhUSEoTi
/gflD7+r4j+md73RhxudA8clwRq4Qe5+hgGUAawYQqpcUCxXzmDuanPN72xgZpZicoQ2h/ASg1gN
v40IBF7NyXS6LdpM8EUmt1ndJlnzvxec4P2CkXVHMmGwppGVgLm27pJg+ZI4URZMHO5z5Z63dy2j
vriWUtPmYaaGUtoP13ImC1pwtq3iC4wZGul4mOGzsUm8O9GqKtHwsSnxLCplYyyrP80kFskkY6AC
SGrts82UtZFv4Tm1HBDr+QcUDpBG6B2ppvUnZY1IQr5ey2a9RBkgbK7QII/M/NnxgnPUMlrLbqVr
4m6L79dWUaH+moCvqsuvMrC5hD5AVhm3VvUXe/YHVcmygeyBooxK6Ax+JpN3K5/dAWnlvsWndC2Q
fz+DSteRwhWEtbkzYt4FsuoA0a809+GAoR6uXnYe6KJ+Pgxjv8Q77oEgJ1SUBgButvB06D6052gA
653EzjOavyrcWRxpvlmxHhKNlJNgHWMkxIVxGsSr2tAi9gVG2pRznfCOypYUgatuZzG9f9kfc8/l
BiKhHDirEvZsQzMcobN1D8CGpDN9RVpKk3tf/Je6uVXXRwqTlVS2ctpXLt8r661Q4QKF76zAo49y
cuABoD126DaNv8dUzUGqAIVAA6T9CRQsXs6O2uroW4uny8hO0DIyPW6yLdSDluRsKlvZdo6OAaua
YCGCeBRakOeRgRVKEY5mtVDT3NmZADA1GwfVBPzudlvqtkYWmVpMq8MyK3zlR8R7lOFEIuaW/4S6
FJAI0hzLuqW0quntSt4K9aF8Cdw38w8DVUXH7nB2xkYh9SQ7sQzz2lUnPt3dv/OgS9ef8FH3WUeE
bEURPkkmr1fInT4kq7pPZ+KoRhSoancvHM+BgMYvTRjPBZfasBCbp8f+TsR7DYlL8gyzc3zmxqzE
IxSo3iLU8+DnNurQC0itN0q03djGXFQODCxHi4OIgRVnH9hjDrwGqR+UPASwhdhDI/qaNX39D7HH
xY2uydP74SYqbvxtJaN2PvrgpaZbbAkGp2S43JpQ9WsNrA70450W+4onJTnOnd30FNOwlFrvNWFN
VXBOAwOVFr/1cdLBN87q+FqZhrX8FMpvSrEPY6bOml+Vbl/jYaIcdAYpv9ENUw8qqsud0YW/tpHg
wmMqLjJMjWp3ReD0XZ/GV6F/AiIr6fEB9ZyJnXNKmpp//E61HD9miMwOpiszidJGC5y4i/qlu6EG
0w6h3QAN8YAiB4wuowWnceCr+4nP+NAU4NRa51i1+faSiJP1lYPlCKAviZHJCVSWIOB1Mra5Qmxh
cKDHT9sJ+BiU9mK4ptGSHud4Ox8sf2UsHOnCe/jJBgag3IMZUwIezOqSiQKqgOSUPWPDfU1QMDY4
ShwsqdevNQwVxXKaJpo4LUH7e2RHnVC7FDrWoMz8T7OU/wP4U71Kgs5AgzgncDCeS/BAlvMK28zL
E2iZ4+dNP4AQpAOjiobBc4QxvH4OwHzsuqqNMlLeT78S0JpDNjJvooto5DMsEY668RhzgSYqgn49
5ov66YPm9X8GN++fAmM8SC00BNokxr0B8Dp93ok7w7PZ4D+kVzfqIVqW1QfXu+ZF5tyFQq6qv6jY
F8dZjOMJNI/IktLTpZbJbXtzXprmD4JQJhPAfy559BVHLfWwG6pJxTJFMsW32QkCVA5pNMJbM7oq
hIFna3ZPPGaNNXQeO4bK2mjIj9ihP00MT1CC8RhoHoDE3klCiOwuMJgBvUnEzC3Ax0j4I3nig4uk
FJmMWO+n2o9M30OIgXzn73ocQZcpslHzXep7DKUErkgmU2mqWn7LS7Fk5qoLYSvy/oV9Wvx+N/xp
XsPEZyT7HBcch0q51qffz7m3uGoF2oJJuC6oxxD/6wM6RDfV1zY8zslrRLO1HUh4Li27eyNCVIRI
BprwZUJIG832EpBhC/aLFuzFcIdztPn2ETm3viW/vvIQBC+CBYc4grkNOTMwv1mqWljF5hKf+3ze
srqlmnwF3CSMMoW22dYewddDuGxlRPjrvYiapQRxInziUxunDKMHeWaMgdgZsww8DrdUQwlIUx6I
a8PXWXvkKLdncGMeTyiGmKz+nUnQQAzrMdPNATabYV0nQDgKb2RGPGBFIvSBZIrrIF/o93PbOglX
K3o3GTMHqhQXMQ72LIzdjS98xHED5j1PFUIXtCeGCCsLxy+eRk8EsjLownQlN6VVaSyIFmO6byZ8
q6KlnliRL4Jb+hRASrZQJptkmN1VIhcZUGZQVqMpycWBHLMZ4wJVrdokdjmTAUmfgy75VU705586
fhNq5sbkoIBTs31KWKO4uNRtKMqtl5CmIvkobDH8I6342M6HFLrw+E8hfPP23NaQsH6+cgxCeSzZ
yxV2sU6ZF4WmH//LnTuSDLhdHHn8twHkYBrcCtU7CtY6vh9mtvAB1J9/DJcQzqPBm21gktCbMUqU
/ZRulxxdK5zBLZ9oMB8/exGq+DHIwN9sRbk04AgGayne5lRIrndGtMq8eXlkYoJSCMbfdjU6LUoA
U/rXThoCWr0DUJnPXoTbZle+pSYChGZ6+wH8B1LIfVuYfCdBLFMyG8BRIEeS3a2bSlGLxOh9MLpg
suZ5erQXYIqrgBv82FdeLIaxN/1jtN326wnZoGMzCZqmPP0efpGwUnSrvkRhT7btensr+qm1oBED
7dwVp1K0wTMEPbATYK0rwJ46DYustcTI6vRIvCQwEDy6+CIWht+SBFDaq6ZybTyJ58hTAA59xgXm
58FlQpTLgJskq2OS9JqwYWm9SkEsMFguJF0Y5Uee8mU04o6sCuZxcpn7nbxRV6Ji5mmzfSublFCm
P2nZnx9P0E9zitCOaUOqvRPM4EHZu+dExCWw1SRtLtYY/GIryUWKwQyK14zq0wF8S6OQoO2uMH3f
3dJxYZlp78L8mog1c9Sf6cS2hPyzvQnI01lLP4y6wIF9RvQv0T1WsnYnw7nKp8gip9OxH2x1DEMC
8txUs/mgyck9vT6VgT7WIqOzF6N5+joyv+D1QVZuJKwxwt3b7iLryM1bKQuwFOksxz4PjyPKYFhV
z5gKPnObhm8RYgA5Lj8WwGgedgY5wIKpuek50WKii2xfTA5X6W6gutNu4aDPIyYzIaolpWlB/u1U
o6ArMWEXupB8wdjALDJCPey9CtBv01fm9AbS9lDyKJfrSlO8ntofVX7+l08TV4oVnaUmkJqVhYfV
hNOosHimNBN8C3gpNKytFjp6LuCMtDnbawR7IltQfwAkfuuRcgmUalxz7V2qXp2Ppx5D/06Od6mP
o5ylvB0tFr7oht1IoEkMbEK8n/SAq5RO+/janfJ8KuZOHb6lolKPojaTyL107jW2m9M2eRHGTLJD
vzGxzxyaTboVCwdjx1IbjNY5TYoitvzTV/b7k03nb+JYs3IQs0R4hdEthzf5D0jnGc+RmqSFpA6t
Lgx3s/21xD1q6s7LQbWCN1qcJvIaUJ7ANGAx40JQyUL6zFkltPK/ICBdvAWuqUOL73wXSBQ5fD9f
QEa4gz/XoFi5TeTpC/iA3XeTYlcAod9Z+4MFuU4wfOJFMy19zh1/ZS4kJWBj4l1OK8wpY6U8kNGS
3KlIGumSy5mg/ZrcsVPAMXwRYBFnZ51AYg076xVm9MwId9Zx2qa05Ibl0UiTpmOh6CF5XqHFbcKs
hFgIOhBN0XaxR5oS2r3hiwi8JsRp9xKKVR3GaJLk3TjGORHSmJ937MoB41uGhZtroYkXVM4h3P9Y
P/vJPOhmuREHO4+oh1En9ZOOnRoid4Fk72JLfOK+Y82zOdjdEOhl46GFAX+vweupn5ecaShEuLQo
ItQ4LDCb5uX7FxjhVwV1OdI3/j+e3I6y/bD3yKJ425BOrJc6LtSmFBcDCf9tUA8usn44fFGP0Yk9
aG5OK/gkysqqsjdGSgP6deO5fXHy7SJmxOCjpJw+mJmgGZF9Oxdubfb/U1kL+LgtLTWxcZyGA+bY
vvrd6lV2ELy6uCqv5P9tkSUXmYR84bWfwPuq/sZBkL0ZUO1zI1T/iDnV2oBayFjWhsHXwSFPECsG
xd29Bpfp1SnQUd5DfbZs8KSpriDywiFe6DUO42TBUyW334RHjRVEWV1s56wiCRNLHVgWa/qJokgN
bdMXjVdDHnlAg4eE/in2Ds18jKFXvUtQMr3z3t6RaJixwljpduaXA7s+kqKV7GQUwzfDoEdyxYqw
LY8mECZMm3+QmgEhw9e5kCdPKmsfUXEzGm8kGEfyfu2rxq/C3iEE3o7ZlMI3YvbLNGLfGqyguTm+
WmfMsM1Oeorhz3AOb7MFt5P5QwhxCs1trh+X/RbuBNt9YFRRG3NfTytnmAi7txONbRMuhTiueNjY
txrUarPIjx0Qh+x0ViRlti8N/t/Ugfcc7mlhFVgcNba4hiZSk80TJ/CvUxFENSRnRAbAc8B052mo
uG6niC+1YGcu6pdXceLBV+iQmeVIpsouyZIB6yZpOTFnmJigbwxRWxJHVrMjNcslptGiXrxWLP+h
MC/Ubi93+9whEPRgT7sSQ9n6Ecd7mgfRV8DMerp+AEHjIFaRVAsCDyscK22eCL6l1qmuelbJBAjR
vQ2GZwUdIJQsVAhbR0At1ry5y4ZMlWXEB3NH+lZqr8xMjH2d8IfNKTmcTH8cTqABvcOfHiSmkuIK
K6z6GMU6m1eWnX5sWaAQ3DvUim2as+60fb9rCj4uZ7dqrHqVfEySYIX+WvNrojGy5jCSrZlGGEXn
vzltqvWwni5oZHablWqGBuHm4q63qewZlPk5muF1poYM0oETB9bPM/nr32PsxvVZl2Tqq3AcPi05
hnRgAdsD1ZE7/hPVDNFuujTJeA+Xvg8ka/AlsjK6ku543k0W/5U5FDiCbP5IUqbEmv3Av/4B5Lp7
gGHmGEj2KiG+IdIbgphG6jRYvJfH0xGcFzOUtGlKu8kvXQ2GlzPLLDGPtos7NDQsa9d4HxlXF4IA
JSk6etFwjOP4Gwpd+kgmVwdU8Rk5X9wwcMLVvfg8TfN94qRYOr4cKujlFD6IpZJ43IY80HgCcZu1
tyg1Eoaav1Hg/o2o9LfvwxHAKKWlvmV6LWDGRGw9IW5jwyVwJR3ZaTSjBhVelYKIaupgKt/UG9lh
AfqOm4DHgAvGnGAQ0Jn/1OPcUJaP0v/CyPJZv1HNe7HCSKfKkkXt4XBPJdWCAi0mN+Gh1qL3Ejwn
tEU6fb95J3ClCsl+kkcOPTopVzQfdZvS3oYpl27Hs8Efx/phGXUq8b6JTaXRYGocC97vJI5OMloH
9sn2F8BC9TBEYvFXiv5gMI8+U/FVsdrQwrNCpbM54wbjdwM4vsBXT4GCr/j0BgsqySjlL21pmvkH
jWCiOJU/bkX6qGHybdpVbSyTF6BJSplkJLKgb8gJEF1OzjWXlxgbV2bQStQL9P7EPs3VA6WcocG5
rGL2GJBeAE1dqgl4FkqTRmWpyuGXkr4wcG+25MkB8TQ1xGktnSMIKMPb0WVlEEZfMeyctI8trtM3
ifOA9UDNcapwI9vVzl/5qJ1ZRN7DRlCi5H9GU+FZW+ZKZWbRPW7tc0XHcTMyw3Yqbb9HTX9zQkdn
7x8JcVxYIuULeMvHn6Hq6q7g4CEpPqbxs8NvgYnUQ0aJPR5r9Mf5XXIJ5ozTbUEao88+5dIuOqbE
Hl2mvzf3uVb/f4yz4hNoj1OVL2iYOBGalfLjR/g+u5ChymwyvrlbmF8KyOjYUebplcUokykzIH7Z
WHV3NXclN1cjuOf+vPZo2Db6LB1vN+DbDdU5mCpvJ8cmvD5TFuabsfXZdEfXQaojc5M7ePdthQgm
roc94OS0S2glqfv9FZ+S6Z0l5A9h32pb4iwjfZ9cF31ZrkrB4fhJH5UPVuYsUloW/NYWTG0ep3kJ
v/xX+oJFzpQy1xEt4jj2WWDOnRENrAiULujKrQIIezP+z5AW1vqgWYRAEAR9KurSsX6bL64Ks5k2
soc7vACtYklnnHgcT4o0WwEnHFXywEBDnh5CB2USyBGjXzxkZNgtsb6/yjhVxXzA10knlx4FdN4x
c0q9mQ0BgLX7WVROsNyRpTHErUen8bHqDw+CfYHeF+rojhZGZ8M4dPpFxkXaGAVG1uDuNXvsIOGy
bOjJ/ZJXjbKbX+ed9gMuc/oPNYQORpWlN33Lst3UOOsp2Lp5o+7n5LiPmP7tw0J8/ZxALduC0O15
MdvuC5XTKgIe44TM/JzGUTASlOb/aP6tq+hm1FE5Pe44CR0KWkDynJ4mSmGo9l1x+uvMViseKbIC
tq5xKndCunF5XSDJjPH8yfDhC4j1F0+brjm9mbesbitqZfnuS4fSAy6YOioLKFpjlVEuNSaOeHTk
2Le2ZkHMchpb/rjNWACyAIyKRTSVuNx9MTfo85wvkvnfkgXVIKAyjPHRca695xY1Kfmfh/CBBnSd
fQQ+lmChyqykZcOtavJXXaE2oZAZP5S3mwAsoCEHxkAV/tPyDatWPbqrLkXeDpEYu0Sob/UNZB/j
/dS9qs9XhINeeuLCrOEAUyoxOSnmLQynCJCvGqvtoKMgPH+JluhrEEOiOcmd6zFFKixpaF+QaJPa
x7NoZrTdTTjYRFPU059eNQELvJDF1aPYR83PYWd+5kUm3tb7ql1gqHcESBz4q1juEtT1pn1d4H55
N2y84hRJpSxM4y8oeW4lPUwaC6ryvai3LIpu5mIsKWKboF/IrW+6Y8zengGMMe7k2VC6aTC4Y3aS
HVv0KSY6/HPHqpNbHfAeGRqzRXfhI55bkoa9z7kQy8UmVX5T/cwGW7wafsw7GCfzhih8quHG5GYn
/ZkRLrzJZFxD4VREPKkolDQL15RhlKs2ZIyaTs21JSo7z4AelrZKplXAT28TWNuhRenH+lF6hT8U
YViNhXKs9HPNvH6B2lZIn8UyzWIE7uFHFO21d9WFEUyEyzD9NPapbmGoDLJdOFNcDE7FersP9Jur
3UKn9JJBJOqjyUpdDraqBECtC4KQMS7fGsTeHyoAb9NSiOByYo/NhmTC7Jei2ShhRhx3/EDyTl/8
6Ge9jPpcI/IVXGTczWYEG25H0CppueE5ezdFGDK7lJUvtLykMYp8IVtjoBUPgIf17wXE/nT3scIA
H3CBfPX39HjrDyLB6kA0VgIRRlB3OnGgSgzhGgPZ2t4Kq/g+UYdQHJQf8ZZD0wnSA9m381Bqxr1H
vQO6c7KfTeSeDijyv6JWlcSXq2/O1BXDzEl4CPrzD038XqwGwcv+vfyI6wAdUgOrxiUnSz+4s0HO
l9ZW66fc8ACPQIDRdPJGCmD36KDLziSvAb2i/PmvllycfSKFqW71biZ54h+5Z7wN6MBnmc9lpyHO
S5BLSpj9TCwJBvt9oAw5GntM1D6UA/9Vl7F8p5xaZg4hFqkDu1gRvaU4kUn/ABVWzPSrelNF0wQ6
Cw7XvHb21uS6LtPZBkh21pNl6iMCcq4weALFZasjhGcSNLuN3ixLDgtzMfqF0BcbMlIbSb0Tle1t
WOswOOSWhElJcWx2qojdl/WMxhCUYFaIjus8Eb7PQr8yL5oIKWfVDLcTqLiZ6W2dxQ+WR2PRHXBx
Bk8BNvcbRjPENhpriDwttbGwvxv6ubzTLlYRUEb53xonlGK1EBsF+k/zVJmhIOM/0ou4Zk4ESW+f
5BOjQMgWTTt1DDfE6wFCrcfajoOsbab6M/I2sGqIuXFwPvI2kRcv0BrvWqZaV91iONGq7p9mPU1V
JiUrRhm4c0EIm1nCyhWho8Yaxwnrg5+kyyUGXO8FG6mGYCW1QcrQ4WzivxbufOhOWagcvgTiwIVr
V3DlJuVzEpSUBS3broozd7nJ+BZd3By/TuKvr5wvv3FzitmosAJuVNl4hpkdNB2DjLBqOuugGzDF
FWZuk0BSyoj0feuEMIw74ZEWCT8Pe9fS5x+6fv6f6Ss4boEJ9n6lA5Qu5gN416D/WebKBv05SHcn
D1AbUOpWVsXY1w6FDd+z5G07SUmjauBDxDz7CgRazhoG6/F+bnberhJTfJB70gAJGmFbFVBZF9zy
efNB2LFPaUHcP1LEq4bZdIWxiG8l05Id9nkl4ECGhah0Wv9IrZEp6yXDy83lXdXtyMPAKxzXCP1H
11Ij1hXMp9iUvA4xMaXS3+57KJQXHVbP4twXZJJPI9XdhcO4rrT81QflRoHscPnIp1k2NS/rvJG2
u140plPAxFgfMXRwsXeYEZDqjKK1AK6rtUhQSnUbpcrAfe0KgRAjPzDyV6S1Y9X7WmFJyOGzpD2W
LTk+Byk0YwtjtcpISkQFEIZNRw7AAdvsOs6hHsa4nI2r/TAl3i4qsXlMLt9EwV27bpDBB0i8iMLf
JdAEERmYzTDYFPWPR2az4oC5umXBfjI9j1sjKDirv5FoYNs8BmhykS8BkQSUKNQ7oxbq3z4zo+Ys
SZWRGU0uZZwYx2uQpqGpAA8vByWl8pVvrZwcbNJwHQZxPVWO4SnHs/J+eR9fxTEu+rOvTW0414FJ
2nB3EfJlkKOKENdPL3QCo8nH25zBnkjf7YZJWYzwdF879OHhEzI21XHh9d1P2bWVg7Q9z5Brs0Jj
AcZYPm3b9+zG9r4SLEyXwL7cSYFnJ9vmrBVQRfTlypF1og99JvC44N1HUC/08h56/EbuZYEcXcv1
gcuf5Hrdu0rcPxToDOejIyKEco373tK/I7pJXTM84iPjrhm2mdAwuBtgEzVJi53sUVePHIhx8JOF
4j32i0cT+VL09BqepBQnLXRnX9PsK837ZKi2zbYOoQa5Qg9inHKbyYB72GFPfEemW7MIILMlueRF
r0P3V96zc1ZQBQNn7VennvS4H+5bGMf5l3gJucqO58RP5MN0f4zbFMkBUfSq3C2mq+9o3aoRlCDY
ymCbxtO7JAv280+z5MTzFEUqp+XmxxS/zA/mmWF7yC6yQ5kKOfKUBheOUYnvVGXN4iQiZzNjhCnm
wQfPr7TilRzQcdWnG7KmFmppqQJ1hrvVMwnR1tLF+Kh7ACAFPQb0fcKCd3cpAlAuAuG7RmHylrAZ
1Z1lObNew8WirGnEd2JB9Tn2sAYsZQEk+mQmkp3d3VA0PIhy4WMIIFC0geMjCsISEdKXaVcC1tK9
ljiOStvapKVmRWBIIBCsgH99ngo17w/rflXIyPDo9H8RrCGradDJXIgvdomTr+Qz8teBVytIj4s3
CjlBaAOWyqj4IhEd5L+EIuJEMVUzRePpL5sgCjwx84CFUY+Ze0EElTOSoEYR+flfKkaC0uvH3sYv
JSgqD8/mvDj3PVykaHAqzQrhvSOlk4soGF6UzkUjS3HVNBFCcvQ6vkq3yRHcjyppJyIME2BC3wJL
TRPBsaBQs1LTg7Ov+y+enrWOKDzICOWMo+BD1UEqvLOyqHlNbWGW+TViQ6B+Em5vOw8tlqg2p8Tl
hdieL+NE8LUp7CxajyIc9jQdc8EMzcnOF/KMZLOcIQGBsQxWTU2pIbUG6TvE0xfAWPkpOsY99Hjc
/3UmyCwJtF1VBsMeyFUTf/qxK0vBcSzIYQxJ3wfsdEFploTwEDszKKCvqCan3fMQ1tPFgUj5lsPC
ajAmozmngG4FwNz5iU/yRVDR0wpM8ZlGQYiDPWYYqBgyHd03DM747f56Vcc3cn1jsHkRhkWmE3kU
5rqmAxMkmcngHK2O/j/eI3hV29mH5cHS/1pn6DHFLXFoT2H9DGg2t7hSzlX/wAgxXrQSRGOwR5d5
l39alnbzGAS7XPSFk298sB6jwG5ZFKjeqkL0T71Bp+2QlTTfKCqfuxe/WA7in/sZW6Wcm/Tm7XF5
Y1ejIT99yAT+Kj26lpZv2g42+MOXrHJBhQpP5DldfChKy8arES0CsoAvcqutb3uZvZiyrFKxi72X
PF/XVKD4R57fD3/ox8kQcYEIkTbkAUak7cergEk3iiLbK5yGBVoc3ahQ3YHGzqgqlVpZuXsMwi1w
0RLUiwoXR197hM6p0KjdLYpA3PzXxhDvGEXWSrllYqyX9PQ2cQNzqZCBXx261UEa7l8fuaizBXtQ
rC/s7xi8dP8HbPwU0UJM2RI7Atp/ZN3lLQEsOVFZUvScOPWKNGOAiuPcaoktiR5YMGGfJa8beMtO
ciJmK7Q=
`protect end_protected
