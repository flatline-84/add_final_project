// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ylOfVfFYyFPW71+laU0Zq+2EpIUc0frgyK7b9byNdqQsBjR1rOA5GLsUyLZjx0B/auw0Tb67ew8J
UXANMKKLJPwyj1u0svPmh133ZU9IckxuspKve5lf8p9W8ptFB4AMJHljgLrz1n9KzIrJtmgaS29X
CjuP9vzdDqZsC7sL6tYlbeSvJn9CgM1tNHIUoIVxBwBy2rbAR9WmMWlcBA+MaXN5aeM9xqG4/e5j
a3h8m0g9NO/flG5xJj9rhHE/PyDMB4uYi2rK3fySo0XRs0f6lRPoxcz1U1vy2bVKWzcCYr+ejDLC
JCEeXzzwx72rbaMQLSZbEi+j7gcIMkJp76A/wA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11120)
YfsZZIBXkGtG226awqUdpTjCnOOdioJnYCgwRFUURmPbPTef0/5q7asLQrl1UHv0BNVBhP/a4kpq
4bwT48jPIF50FWHyyK2jMNsrlS1wntwVM5Hw9CS2kHoqFWoUlW4ZFPOz673CvP1o71FZvBqcB//Y
OXZNo7RXCFQGUMNyfy8ANRFZkoyFgWqBNjQjhvvMnLs2FWGtT3NEoTdXho0kgnmGe2CbJnFqu0x6
OO8DdQC1O3JPdngpImDwYhjzul5qliQLhjEsbfwNtJHi2ViUIV39Vouevdu1PrVrvvSKj82gJ9ym
I0P1rolG8FKoFCsTw9jO4RYt8Py6xaEpELuTFaNoaiN2xnS/msVgfY1OUKSSBHIvwaIcAh+b5bsZ
vmAbkQb80N7f7jZ2B/rXvz600QSzNen1Sd+D8b8H8N4lMRgDEWpKBlEkFXLgyplzBvY6SPilQ68C
UT/zcY2vEaRT1Wnh+0kKgdcTTf5xIJxZJC7dFuzY9FOKS+9r2UwhfnuonPdy6qBagFYv/wkTljW0
ZHPrhiYALDwQj1GlDimhLufPdjYlUOejI/WLr/95iuj87jCHQSTcuZJbFaJMZTt9WAfpzHVfvBHZ
O5WyGGz6nyMocluo02gbGKZP0pt/7xxGZ/9jICJiQszKpD4fQCu/xTPj90juTWPuf6ZePeLALjzF
7xnzPTstsxIf77wmH/Q9zjZNYgmmP7/c5UePc4bXXys4wFd10zA3LLfxbryr4Wu5uX8uXJXZzgmB
3xjM95TFnz8a2YvgjaDGk/fhimW221bpKUx7g+yUUznv7cB+PWIWqRpxlv7b452Ll40LyFtGjCVf
q31uHCINjV8i+TBGbg5USC3iaxKVtVauCqt0DOsiWHu4lO7N0nD9wV1x9wEyB/NfhlAvTt77uo/E
7SJLJ8yhlgs3w7VkRywa2BAkcVMdUVIZj05U4++FponbTCELAJinvx03+st28ANOWlIydBYfPtxP
BZHXq4QdoTRbLMCLtTODDU+UB7KUoBbZks1cRtvmtc64oK3oi4adRmbMfklBZDtQSWAaNhoFZ2LJ
penA/4YtQ0vNZ7sP4acp01uLfqkoFUyxrX9L9sQ0LuheK9B059JYQuSWsaHfmjP2foz9/0nCkhtT
sIRwJ3hwphVXka5yUo5ZQNEq2PXKfCL5wCMc1A2/f7fTy0Ib1fNkwF1GBMe36MB1ugYIra4Tjsb4
P9yS6d+yk6zdLs5b4+HBXog8jdHMiCo9qbxjIuyKbmouNL7kASdX6oWlT7mjdI60W87U5sjlOobv
G5hFSxA+KKRUC6zWcwMBfdJqD1WD4BCFvM7ehWmgqBDaBs4NEnGUaCPNslOVdCQRgz+62+NXcKwf
J7Sa0VxrFxqbWqIC2zfltb/lireJCQL/IOiXsqQYkm2Nr/4bH9zZEbyKTEqIMkz1USIDoHnzgKFL
cp5Bm6viBLXVqZNvSqkMK/fmthB74TZ9JUpKBhSomt+LdyW1mA0aiBW8XFKJJKT7yR4gUOjTvCMj
jO8FMGatqN7+jDSYJyny4IblMNZbvTmNiflmnXfN/n3mkdXFkEE7CHtNCNYPZE8iNHtNDDfzVio9
nFb2bbN4zzgEyds+9Q1eNU8M+OtWiE8kxB9NVCQG6iFpGQIrITazAGm7+PKpmJcHefuufkuJXD+e
FZaFpFPi28vcOAohPOt8TYCW0fbyEHI0/kdURgHkNqY1tseQ/J2itnSdTeR/7yrPTwofjCBzi+Xs
YmXCsTBNjvo10zj3YpEPfel/SsE+gnNBqe72hj6JVGXqFzUzntlT6mTu+XF+UZifQnK7BV/XyK/E
/wvF6mNx7RWmZ8QwMdGezbt/Y1ziNsniJuY2aU/e+NTtZqvtzMIVCWR2vjlN3a5CqYJwt0sk6saw
pd5QPDyKnUoSdtCEH5Sp3wLmkQvaFK9blW8a+TsAEvAwZ4B8zwwa8HYgmSocm9Ufcb2XFQC0aFQV
xf/B8Cks4jvyFmCnu8y3mS/P3Biv2WCyprW3NhOnjMNJ+ddoyIWuK5/hTJK8pbSEpEXideMD87M6
IM5W2Z78o7965Kw489RF6yR9880qWlt6sEwpo2erPymDlqsPbLQw/pxJHsSDGUhWn77ErqVzJbD9
v0PqHpNmSdrr8vG48uiEjHvHdPPy/CmQvAJ2u+RhVICKAj0PNTC1RLQTLgvrUfA/bc4lzQENacb7
8qgmIhtNRocgfzouKkfIj1EzqgVHosPx/NOKuexoiSMcRSFzh8c9oWadykayAW6sMGHg0mlDkHrZ
gWAtOBbJDJvuFheplfk0DaLZZgsj3HK+OKcj8M90+DFTH+o4AAaU1xICdIwxqH3BZEZozhVxifQ5
YvhycQhk1Htfb3bNeIWF5ovqItj1r/suDpwAcAQYSDEIYOiTuUQtU7isqM5ZGfpZjrbLsQHlE/ZT
2RfWmDyvfiXUfq9BFybYgyfKlXWT2QPfG4iDAtaoi4jcX525b3iVbf2n0fsLmk7RXbs2vWkiDRtG
vBXu9U694gIYAn9OsT4UTDcGy87Qr8Z3tEPbQ945I1p9bcC3Pb2ghLuwQZFg8RAIXaPak5zMaNsz
JIFfTZNq2JZ1mBRPZUGaS8C9DbJ6wh6WSrT2cSF3I29RYBpHC+RX6GXDoOX4zO3jC1TwGfA9lK3s
Cy507DRwUiYixX+9gpsfitLGEK0FykK2oAi4/T5i6npG3cd0yZ4JRCAVf0h+qOKHraiPpG65b1qk
GF242RHq8rNNdlKyaMl8tDJRE07+dZ8e1QvK/aAnalUZgFDAWNR0LY3NXzTkxFeZqtLhtosn/SPm
B7MTzqsDFbY9KOfXDWKxehnjQ4AVg7QfBMiVFjr3s5gnPtr6Vv0WUymNO16mGGg84IcK8KwB7Rgo
gVJcUKopN5X1fuXm7O2gWU/sJ4RGD25DXUC9B3Vn5LUHENhrGZTzYXoTrnMLPoKnx/64HRiT/OX6
OMyKQrD1f8QwyHjEo64dYt0i7lrTWHBGUa1aovZmRQ2ARjHKg72Q9zuk5OWh7dqBB9ZOFARAN9f6
4zoG1ZnYcfJBXOqSTK7ixhoSGQtEqHoDMLcygaybvlA/r8Pd+dL34EefxA/wR6TDFRtDfxRcS6dH
HtFcIUoV0hD0hfA7CClm028ZoLMUuz0ZxiYU+u/yda7Eyv+jXEtqeo4yCH7wx3XTGayez5EDNII6
GPWqZBOMvlRu4IXx8Vvxhnmura2VhxISUq+Nw1rx779c2FG70hW4qF2AM6O02R+2D2JNL9urSZVh
yj3aFpKYmbOt7zH0t7EPkzEADpSJzZrzxsRwD5ja7dWdccNRgHkFJpgpXr6Xye9oNUfSZ0zrqcvF
k44imsL6I63vz93XxPMtfbDRItukYxrJM5dpMd2RzNIxHHR62lGnyCC2pH5+kyt3TyzNdI0/uYPp
bVEow1Hwe0J8U1cnmYf+GETIqAN19L6t4J4LjRaMKrnHEXhLfUHRrwVH3N9xl6KMA0CGKaMe8reL
tgk3RjOyjHwzMOjsmIRjAzdQJHWFTf1FCXgEf4XJQI/raD1U23lsK437Q97BqwsgsVd0oHse/JUp
0WGJ21NWoMw+uh2cgxUjW4gO9T4qBGvaDeBlws0R95N6m6LhzNg8HatDSpWCPY4n3KIHBzuYnISX
oMnTBrl2Ey/4tYGWohp4flVPxru+e7RXIqtr3HXg8AYzRuxGGYzrgos9g+FZbtxoteo29yWGu/Iq
xXuamZ+pUcQOvld5b6tBd4YQHXjT7ow9/nb/Wn/FhyLJAHKOpVloybLmXWa0Lh1m3TEAfY1RArGW
WMlNBPxh7Qs/ERVO5yyWLXK19X2R/YgqWK85197vTGIVy0P6ulwJ5Yowx9aF/J8j4fOdWYJ+6mNd
azDy+f9zY06KdzunMNJbcq0Lhj0US+5mqXjOJOp+yUwzGrrYpjbH6LofAf5vXcuOVd7Be/vXkI/b
tDWJgDrkNwwRnCsyhb/ZwfaDGs+pAs/chxi/S4dDpg8PPY+YMZZOAUO8dKH+ibvkdoOT/GxJ0geQ
8nWP/yPvyobFXUYCe4qd6VS4fbCGDo7XmpwI6pZghdGg1B9grjulGvJJiJPsl1RfEBMgtmM2jiqU
01+3RhENmtipVjpAQD10m9Wxt/oYXaHFI9ARM4Mljgcn2aROXgCL91ae3SyPqyw/SXSKSahMplUf
jfzg1MzOR8aEw5k+d/fDtK1n4khj4pJ5wfqBKW6JR19z/rl/5V+QXwFBntkibHdwrFpIfeSk6b5i
EMO+eSfWuUuWIGhPTgCQPufAQvnfc5vpXjtU3qJWZoKAkwZT00gi7//Z2M40Ra9SNlcHt8xVwykY
dKp8UsVXJcihF/QI87jZwz5uYG2diEIX0ZF18ku+PJMpOpNkoOVyxUUQIHuOkyAfCcfNVaSAbSk2
64eLFgCFAHGSEdOflj0RKDQJXAnypfyOUQ9ENDh5iOvQq7PqyzoXAaptXZPDN8vzBgtrJSH1PueV
SPQzAO7hAzAPMw0p7gi8Errb6c5gqDSDlrj8YaqeSXVyA8nog8NqJgBrd7T1+VA9S+eDIU1nkUgT
coThX4wieJLPgLZLgiU1WCGY24KaxFgPOvlcvfhpt1o0gKZHRE9RStNA3FWaUbW8MQx4Xl0fXuJK
09NF29rWbrg4DjeURjPyf8lInDRFjpgIK+M5J7iGX/FmVRFJ9SclVpsN8+HvOs93SvaagW5yi4N2
u81rqIhxSQsM86nKqKf7UYsHaDe7OZEwDR3qDVj7x/PyNkcFefzskDABtcT1NnR9mrjl/9dIIbAP
G7gbbRWFPuzaAiVIjW3rBIpSg4Gx3EAH7BVjLAFgLLQ9UZhPCm6oyD8hC3/BSgOCTYTiNH7FECQI
rilNL1YRu1Xv+S+tg1MisE+XUEsaNvsGMaJGLLe71WW5lOIX6e8VPb8kaoCgFGivvED+v7JNzKrs
JAYC847Sc7Js9vIfs67eRNs146CNyrhDZc+1W/uFVVbJAbp3KGYU/ZovG/pWVBOCYi8O+lsfFHKX
Ngjx6LUqE7PbLLAs0PQ+/52xqfB6E5LfYdRFGaDxPBkw/GFK0bpyiOkJkJ94r/XZWD2b6cIURr58
iCELKJj3YHQV9BY+x8n/sMkqwVTgDCB2SG2yIRkDvfgOVlyidcUs7auzijrHdMn/ACRnp9ugNpgC
w7YpbqrP8CvwSANX5E+fJ8ekO9JS1+NztjosJNGxmuKAo9rfQj86HLhaWy5JkyFBL0yXh4X3q/YE
cOtCxi0gVmfnXoI5IWzMZnZi/0K2HRCcumGTcU6VMmtgvyJkuXx7XNqqEwrA+mUQ/8V4kq8rTfdR
1O8rU8fLCtH8WGUdXtkzTjV6uhpLGyVV5ZfkNUEpd1n8OTI9lpFH0Yyl1u3BWxeugboLMm8CFyqU
J4ehnJDKiIdI9pCc+RU0fHiS9Vlg6MZI2ASXABQKskp9ujK//D5euN4fJNW4I/K8BR4wmrJLsmF6
SK7OjeaTrJuguWa9ee+J2tUapgcuJeGfbfApsDzkuw8vXAr9o9mB+dD/uKHN08wr1Vi6XtFufzhd
2xQCj2YwGOquFu6eKJOIOIPHhRyw2KDu1BthYvGVx44wz8D7OOn4g8G1RF9UXMcVTB6Hs4eKE5ja
R1vEthn8UfEJwxm0b1L2bb7fDnhM3rHiF3xqIGWlt73otFs+EOIDsZDIFLQAVYi9dSkOLJRbUVRP
PWlTMx+5EDo0Gy9oKNIvMqJ5X3LhbBb2l2k7lQ9KyetbgdCvL7BAsvguW7GpbFmSPKOtHE9Mt6Ur
4F21xxEihW1C6caTzPiqU9w9wg1LylNCAUCQnmD6RHvebsWRnzf3V3ge5KhG8Dcs80zhM0s0vmIp
hH0D0UhgW91skeyVjf4yEHd2wj9y0HSuDkqIV0GDxODmZ+0fY335ELTBPHEshqar6PvmM+u8YUfF
49j5c/Is1nlNEmpKdIg84tPQXOagYX4KaGN5GG8ZucMPMeXQJvWt36zwaPZlDpNWcSTcJeYJVNZK
J8510ic14ukl8IGmUt8RI5TO4RqRJnlMqaCZaqph3g5aQWB/dZTq19Qvtf0IED2+JtmtasxZ6mdY
m5EFNfIfxvxs0r+E+ALSQXLn57aWK58SUQjZRZzTFigtu1Ozzk2mR/AtzD5JDQaX0p6lirDi/Ync
ih099DkYpb92Ooru6k0uClX+I8AoXAzf/93QJh0h0D/hSVEBQHPmCRZY1vntzWSN6AqjiWhou5L8
RG1cWgKM9FhzEfl2KHPb5J1p4wXnIWBnyCg5uNbnUirSXlYEg8V/GcyEiehAnsmTexMvRX4N88Ez
Eclc9eR9/x/dRB18y+NDJ3Q9jo/6t+TPhT/2x3+QIgSpENSELyKARKfBCB/IPiAgtqnJoRvlUPI1
kY0fvT4bCmWxCzExa6ca7SOPm+go92DSPU+c8GUNk5QRhANVPXeKu+9FfBHtvmIO+5gNwsHm4dQa
UcFk6VYgeC8udwz+c3TSdVWwK7Jvl4IPezSj9cjrAi0k+Kt8V7N1JrwGqP4CqouI2RdfTHIhgYS8
8l2Tv+bmVq5sjjPdl/2QESLHi2c8O5LCoFIl0pfYljJeFr42Btm6ADNMF22PKtyCYx5mrQTrhbSB
99Y1ghbVntrmq9lStljhR7fdWgDCa27D0PqAOYqwBLQ4E4UR4gPuBuzhcPyIugJ14gs6idpi8aAP
h+CfYQqZoPkG8J2UCZRtvhA499BCCxZBzr4lbWB/ulcodrR10eHKkmmp7HBOWyV8QtaHR1Ob2zy3
dVTJmlUzNGNuMHMw5uHdgaSUiWJKm8smp4PMQSp0hRjWvX6+5EtVutfhh+dpX2fiTjCjlsctOq/5
jPzntLkazDrtOVKx9zU4qeb1FOOZg9MOL6wQfaotTRllSOd6Vhod793LuJJcMDF3MO1oAJzky7/b
U4gQ7SXmfrBafcSOKHIIFCsy5ItFUeGON5eeYMkqeeG0JAun+UI0j5FgGqZ297YGlIbdMkfaDTKH
XwvM2Mp9i3ee9DcNDWnyL2NBsmwlCLqX8jP7rj7jfp1bMtzC0r5BKN/gZ5K0rQMKm6jMxp+28xqq
pG5MB7nS0Bq9jL18hTswSndfwRmGKAh5eJXquD8+xHJEKb9/kB6/XdVzw2roWANf5fW8zFuBhEtG
qV4tBwWrH8478KJdAuJ2NTG3PfW/rcv//07xXxd/VTdWPVyWQQSPWYt6bQjmgaykhJL8vNOWv8Bp
HXLaOkLskhEAJCKT8KPyJ0Nv3tH6YY4XiswuEINvqSujEvEWBZoyIdeZyrXGeAp+51DwMdm0OGiB
E35x7PdWFykFhf1NVg86cZY+YHMRHqo6LwHsSqDmxHNCaQbMEne28ZiVoKhTn1V62ym5K1amWIEv
t9Bu6nCPDqryLhVrapidPJ49a4IPZ69rLc4zMQSUS9Foz7RjWTx4YsdKtotsCw8MAb6WScvtjWY9
Er82P9WtBtxlzEcr8T1iGRhAZbbQmqHtJvbBtUIZsMY2cFyXocGrJfcPEUiduH/lgkBo4VR62TId
w7+gb62ux7SWQtIltK3MFiu0RbTqAHd+jBDvbSnQbL1y6XKJjF5w5aPwka8PF4RhC8xS7ngnRqHr
HlUTMW8mOWBlLQZz+wuWyquGYGLRgn+HQV7uHeQYgzOwH+GDq93VYLfpnjMoI3EyhCeycmJOKsVt
iglsNiIw9lLC54O6epc6yiFgvo2k3VUy7w5FiweS1qm56pUv4V6Z97vpKNcYONCz5Dcj2YyFVcLU
2GXaOhrKh7cUnwHggo81djGZGDO+/YqFXwkNs4LlWSu3EW/9WTPALSROTyPj29EfCD2BWXeXNw56
s4lEtEsk1P01NnphPJYYm9lE+XoIvLsinaL6mWwfSUd8IJV42Rc9Il5vcIpcbf8VeAvSpW/1bB6C
cz9BtqGZiaybZJB4H+JlCXBr9sbJm5Lt93ZU18cP7/NWg2h/XzZR3/Gjf9ImEk3dSbloIfcrloZo
4IaAUFnmzYUG7bGEiYxogCY72VTuEDQIa8uH3SQeipgstzbXqHPcI3PqzI7/cmSxB+K8XZWClWFk
kYS1C59c8/dbfcRNu4tA8jdkI8dAXMyZzAxlDbL5gndbjPHxlTMVUizNyx6s1FJyHo8JvoO0aFHD
ZopkrMWBObgZIrFhy+mg01hDjEDFAMnSShJ3OlNwgF25mf3Fts62Rzz/RIs9Dd6NDoiwSoLT/Oyp
wBTWgwOfK8Ehcm3Ye8si7+rGURTxdJJzOnQYfOSnfRyxGm7RS+w1S2DQcj8qJQm0LaTpoEewJD+4
N/vQ7WrFGpp+mWDLNoyVjGasC5Hi5VxPO20KixIhpsUcLYB8EKfsbHXH2b/4t8rDB/7D63XdSq0B
ETDL/I8O0MVFNzxirX7fVrLTNYSc8nFUjhCeYFgL5KqkjNKKJAFt952ggxDH7VAxj3wxljsl0ikh
AfQfRl+QydSFQd9M7qXjKa7CIgZXf+BmYJkaNHclUGgTy0YK1HcCp1i2WhqxhITfM3VX/whm0QqF
QqlZOG8oU8jQLo2lshA8N1Cas4bBWeNmQfBTM/BMrLCXWkDyOY32/9CwrgFqgsDFtmcup4xjBWV9
ZhaLnlagVQrwa2yG+C/FiRVXxiQxiFm7xPy9CXWeKalDQ5DTGpjpP0ZOAm6FwIVcdZTXjqyAeFQF
N02+opB05BDOS0rQu6COdwT5yOeUtRMrkt2Fs+D2V6T+JuA090erx/n5PR6HScd34hqMXLCja6Bb
IiRcN+y1QPX0NK53iApYpsAbqmYmMnXlX3F3ulDi0rGLoKZfPoofK/g2OyAh2/foMfOSHgY3MOB9
T/EXxchiFsDUwktERVAunuTa1/Ben0lG028xDtRDx+f9MMDingo87fCSPrCBpSlgOsH/PoAG5ScF
KwnyegVsSTzyqjXwgCEm7yBdgKo8E9kvhPwSOb9huwSibTEJHsmXI7CglfYSIgh+9X1GVpJeJa3W
fMt6B2RXYoQhtW6QbRYx01Bt/UoAuAvBrZzQy7A+MrNCeogPbeTSehFJp1QlpSLnJUw5QHDOFb5y
rnhHaMn8ES4CjACWLx7Ln6auFynAYpI911tykgSTM1WVb9fKou8ZC7UlRhNfzYATH8MCbOJaYtg5
Q3U0zG8J62ERBlLfOtCuLzLNeRQPqJrkoMVIZ5SC3mO8+3FHgd/TC9z0zMUW4HkHY7fugpNVMrha
C02sMFvT5EH4Ilvgm0S/hve3LNquHa6bvDXrYUV6ofTCw+NGKL5jgzkwUp5l+UwNVSc86erYNtuY
NS8EsArYrVkerPTXWzQouZJAhsN5B1igTra76NYTRQ/pfIQXzC1LCVoN+Jc4JvwlXMogQy2Jog9N
WDokRx/ckhKdZ3gBiMQOyXET/zOTb6Z3fcBIJaU7w5ToPujI+aiYz5yiXPYcXeZqK/10ch1s6uzY
SfU0AxY48MDLKVvnAg3vyDhjTxcgQpGgJ2LUCWZWLwHnW4PZJB4De3x02mIXBM7aCibuRhnuNmp2
e2FKwNIsTw3h0haC5Qfr9RdmXtZPVB3l9Frbo2+Fnqa7RgGyD/+owu2Uybwnqwdd/aTW2Hgvup/Q
mIAWFSYWQz4FlUbQxdZ9bakTvyvjVo1cqlBNODfE1NdjIbqNZ8dabNNLh3oe9lJkuPCwILuMATXW
KLDOjpC6btr/9qbJFssRfDhgkhj5uaoJ94nlyURoraureMjJvHQLjQOheVKk71heJ2+e1VM1zarw
STZ0G3wazdm+8vKY2XEW/1U4vVkurKnOQiWpQg2HmxJ1wEb+bammfAjHzm1aXfnLyu1YN9g8iyMj
5/dYlaEBlALlPwOQWGmfsntDOpRHCxRMMJdc5GnBgn5xWVS60K/9qN1nAH9GNXLri1UaTbRhxLWq
Ls8v5qeU79CYB3/dAUtFynlWBEtMs4eIWA5KgqNRkOeSNXJsvZsF9wZPfCi1ywd1X5ToM0VTyaX+
DYJ3b9canYnHgkwA+Lfhzu8zjYub/iJHRb/MH75tCgGzu5cOJtEWDqrGdcKUYqJZnNt+b231s2R2
e/uWsRHU36JyKTjCFBuelYclXNfDJrISMazA89yXq3znGfUMDOdHpGAJXHz45R0ufhytHeAuy5xc
03oD5Y4IuiTUp6lvDt8DUYlSceTeTiYQ3//h/9wgeRjS2ZCa62cgLMPbTsEcKdnu6Z6zrTItLwoR
KUVZbDv3Q1uQxGylOhPmx+z3YdgP0a/QAuXYO95liJLJM6H3ycJ8ZAVssbO3pSr83LLbEpLocYrX
VJQNAZihmRSHt/tQT4g6Ep1dvddmpBuaPHVrwf9COywjBCCQZnLTK3AFRIESOUmAYQVfPLksBhW0
V3oNeM0V0pmoS7cs/IInngO0qhw39kCwo3x/cjQD1g/V0/C5lq5QZAtAWwOf08WdRKgjx26Zx9ub
O0DA3JHAqC8DLOmKSEqElPbH335lRHbdM3EQHnliUjsawPDIoL5+pQI3qiwYIniM06H0P5Evf8WA
xMsthEzN6jO0NvuGXJJPG2Rlu21dH1UjNZ4KOLDpAQrL/D8sfp4jLzbZPrzmonuI9pEw8Ut6/7xf
aCQaTwSeQzneYKBEMGfWI1Fv8ZAepJxSkFeXH4ODDJS9iHpoLTunOpYYqEenQ9/Oa/LLrEPdcStB
5ys5+waIl1O48rnXEagusnV9GGX5LrG0QK05DrwDOdLqu9ey7RfD0b+RAMOBW5VW85r3tA6fCUiH
AO4oz3AQoHszIBXaWXqVN2CtmXhCNU7n8M2gBrcMwZQN0lnMp9aAoPumF5cbfSTmbLA1PRAPPWdT
Q08Icd7T6PnyV/xUD9cir/NMqgtKRxAaVELpmKjUJ5UFuCFP1cSfbxUrHS3OraIC2/9k4FHYMVnN
NgeBFlN+Sx7d8BRczblkbHkGk4JZb9Y9phfyWU/mFL3J2x9y/OZgqYaTXpUoxYyaf0j++S/JD3Mc
qMQjqkBDItX7s95E1vB/zNjLGyKbPy2OMZiFumhNB0Ase/Fa3rUtb18SfvjuhBqjEbDBUFOBUOtx
5Oc6iwelcKy6m8AlfcJ8L5XkQhKD+89QgdSyCCpytEUdhHvegRC5wpS77DsR0ZyozfuedrnPS6Zb
YkL2cv60Xfdsjzv726REz3qSFzGoMhJn67StoMM7HAdtBJf63s2qOlL4B2BWy4iCsRkEqLBw+2O8
6DxiKmLKHR7LivKnTGwwjhjhhr7uBW71Ic32xr7FyZ6U6TyWjEmUA5liAKjA2Z6QYO7vL+Tktyc6
1Wb7F6guwJ6gKOkiM7ewXKGFw6l9HH5zavyTHPNp+k6EMNRdHapRkaL+cwG1Q4LwL/ZNuJwV1crk
jBWrz74r/4CO6ju8cvI2JccrDuA1EurH6kXtnnePEcUtnHQJyY/xCuyH27P2d+MbMEfhymT7kJVv
KhbCbK/Snk8gL8CHjZob6N5Vv9lKBAk8SAJB0fnTYhc7G5h0D5xhKurv5cA3DpkVOl7e19y4lwiJ
xw3Igw2rD7KYIIx+bLMUFhJk2YFqiJZ8TAzMp8jUMZ8Ifvg+MEmiOFxTkm2TZ1y/FAk2YYXmHmeP
a7BPG2qMBCVIu7b9GWEVWfcnmS0kcwCY35AP8HFIxhQNPfpM982L8AOuXzhRWA6XUztJct/GgYYT
qU5G5U9TA22W5Mo/zqHRBuCBja8TNmFBwc54kkO7LTIzfLMZAWXFoJOSUkA2FQMLlJkGDM+f+20Y
Tjcv20trTI4OywsINizSXqp6ogVHuP8N+h1UW3MoVQkZbc2GY9GPUB/LuDKUKF+H4diBUwQHyNWp
/30GXpy/pA7+f/1V5t1mrsTiwgejZzyUaO6T5utI6yPodkRn4XDlHbxgdWPeiPIOQhQV4ZQQ0aoK
mmkos3552QTQvrbcZeyiFvJ+m2G3bNICei17qazQ5jAS38jVoz+rD71Nd7UNIag8AV+G2KonbEX/
j9X7F3STmCrt9hqXQTUFnyeUnyU6kEJeW9l7PxM3PztiDyl1AO74TSqpy7BZ164R5/5HUxHIopQW
ndaeHBSiWZU0qyWsckddd9jif41VNpVpHVQMsj7P/LLcJtYSzyLbRroGBBv96ENCwXwYXQTJY4Az
lRwErn372tryvrWCjcgQsALtEVqFHDVgTiff+mzoDpXuSI3JkZD2xgt31CEjmc8U9tiqVCHDZvDQ
75+J/pg2X/RbJqmd5DKDHvAxYSdqqtQOF4KDarCYZFdurSMfZbi+YecuBgnvL7uXQGTIyoWVHa28
T02eLw8YFHjNMTnvd4nKB97HbsTgKODEwNTfvCmuW6R04v1FCz94tWNl17+UmOhYTovViBx11YV2
7aV5e9Zcc8lwl9FxYPBhuOXtBUFEz6ii6WvIuZhch0o4kxCVpX2oZ7gJUUG2Yl1cqSCE+FWYM5rH
usLUyFYC91k6X8qWTGkeulV+j3/5qUdeipwdh9S2wBCI4YJNMm198SIjaPIL7Ap2xC1ukjz2zuys
80QNCRE9v79LgK4JZn8H9ebdJYzP7bIVqriW/K3SdWIsCUChe07emPNjU380X5kTHTXDYGKQ9G0F
WGw7JQuG5YA01HerK4Do8gaeOiDeRG83EqbwylFFYJQXuDUQCEYIrqUptVfkZUIz5LhZqo17iVLa
KOCrupDDbkIvMZjyIPY0hpTpUajNVkTNPfD2evH1WlPkfyM33dwBx2HTAdq68TEmQA9E1k875MSB
j6+l7k32Krpat9JZcLM1z2CtBLg+iAL/35GDHWuqwY0IHpZw3K2n0mV50r+0sj6kp4WxEOjgYDDu
tbuvXsKlbbosj7GyAtlMa2cI1gjQDSmxovkJtiVAqqAzDIa2iLWHpzilgNL6y5yfiq9ajoMpJ21F
OLV8XxfQPfxUMw5e+5I8+zPnBiqXNekuNktkj7nSCd/To+1PZhRNi4CwqBE7EeO0VvE9ZeNusI5f
YDpPCw1cnGmf0tyxMN4JKje3uL3JtEDzJnBtgrWDrjgOs7bVqTbQLfTyvHOAf7v233ThB2u0lbuM
bnvCuAO6ucmXGzxh5uMDkQH27tYTN3lBHYxkF0Dg5+528FwWWu7SMpWYg6XUivVimEbUbIvs9C4o
QHkLMUfvBOreY6QEF2Dgb4wlUezlgPaHEKqUHovCTuIv+XFW1W5uFsJaUaMyiE+vKFNfViCa7rY7
2cUmzQhXdaGVKMJPMny0tNv32c/pNKxgeWaTKKxC7D7TQDU9Uu/Y387ydjRhvkLyZRT7yIHzO7Q8
KiuAf9xOS+wpgU6ds1VlQ5QBZS7ijhAeKsFg9NCoxZD9NhyahK72xeJMvhpLAVw/n5+9a0Jqmtx4
N7zEEVAUxC1uphnL0CYHVtOtHJsWICy77HLE8JArOw3LPLyfFr8rXTf30t3pXGPscGmkXuE+QxPc
JBGoz10HVMGmeM3ciooKzlF9nwyZPVDbHBw1r1VLOt8CgQTD6zVwhyF4hBsDnyvt7xcUiuGtzJif
gxzQwS2vSsAZf40BY8+Wm2jvX9cnFm2HQsQ7sB4BcIYvPVXX0dR3MqEolJC2sAmj8KDqD+JXgBKQ
HHI4WGhOpviOLtWBgEK3xjHQtG12FOBG4hpqxuRtBHh/0Cq2DjIVlZ17hoVLumZ/lD41FUuNLViB
WoNP/XvMg49Mb5YFgFuRXHsjoWUwRBwOlMx6dbMU8YqrtDc55GKlRSA5/yrCAK0sfBrjtb85RQKI
YXn4BMUwn3Fjjf1eWysEBpwcNBAgXBVjXX6YZsv1Jh9BmGsJIt/Trm+ZxujZgRf/+q1Uu6VVynIS
gVk8PlZulHFy3vm7Lgst5pDEVdERmJ3yw/7wFgOFPTF1jbuzMP7acnFDLMzx5M8FXEpq5/wRipbq
r2mYSDlWgzMwrAFM2linOTJ99Ip1YZMv7f2vyywb+l+eaSzv+er1bOoieVBaXFIiSD/5xRpJFT6r
yQk8fM69bVr103OFcVZdJbPMhrtiygxwOVV7WLq3X7A19O1o5PSULVLZamkxDpvdYcVmWgMpxO2g
Pf9SkICefDGbSdqn9DsHnLvGGA26GE61ZftDHT7/crtA+Q83pMe4u/GcWp7OoVyxbILJa+m8XUHX
CEUCejdemtrawVCQ4qhUXDWheKD7c4ksiXvHqLbpc2qpFxM4bmEf8IVlTfxOxP4PMmWNeFffRYiy
V9kagWpReIlNF53qWz9pr1euw3jzC56y7+XAh4PO/NEPiw5rGl15AVO5WwCnXn2lVACAEXa4zCaG
Qc6qzVpYM4D8fhyKZinAqPDZNCAjvXxDVwq+8mtsJkyrdM5zHabXlBrO7j7nPjoa/AgZxJTJgFYA
A8aNkShMORNpdtr9od7qpAal+PePGsTRUfGYKkAk4Wnem1yu7LqDZhhsx86i6xFtbSILO0acWhkp
BZ/cXcNgstwVvr9cX6mgs9PCBl5FEUTd9aTAch/TsUByvb/UX7ropGmUAooz8zL9pdNI8fNRlp97
mtSiA6LTY6UHsF0rfwaVNlO6qbMPXCXXLJtLDsGd7ad66dVS5efFSGE5i7KpbGbl8aPLWfU9BC4l
vcYTWuY2mvolUDHOb0cbQ4S1NCuESIxn3el9kCnw06Sy+9xKS1orAl+hCzivF8X+2/vSCRwzR2v0
mRiyVOQkntbCMCQWi8Uwg+J+oAgsjAmFqYhliL+PGdY/Wm6aFp25eyXf7tROTVfYg9pS5UJRREI0
ORmI2XGQd3sQtYNLQ0/dyghWGvvk5gbGqYQiR/320WRRr7J/SV96RtRrwYXINLji7I6U+sjtI2mP
u0uHlMYO+5zZoC4WqyE4ed5wETEAs9oXAqEH/RKUQ9vlDzU5C5IIR5FVemHyk3Q55HVBI4GZuc2j
t7Jx05Y=
`pragma protect end_protected
