-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SxgwTJKa7Trm5Uz4Ch7wXSAGQAm+Vz0TuSdnZbgYORAh9VJDBrdSO6Aa36J99H5128wmqCrG8cTY
c7CAX83t8R7KICif2+LbyPdZREehhlm0NIi9dQimKMcTlF0plWFT6BDeWNuJSlffWqEZma0gBzSy
6ipZ8dLjGdJ29uFZV8YzyMLCEeduzX+uwbX+lksUfO4hcq3AMWoVmBCTMvVFoVOiZcfDYDyMGxFx
WjBdejdtsYs6F2rlX/SlbBlV6EGixUBAxlNSBKZLlCkwxwdYxzsLJqlFWseRJd9onDt4YfjXiaGy
ksem1FfdX+0tOEcIVaryDDxKxaRTgCbJ5NlNNQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18800)
`protect data_block
ciYyRzuMlJQy3LFnTK3ADh1Q+BDcEqHqHvbRgASRFnEvAxHxSdoN32B/TzgMmzuA2m/B1H51AEeo
IeMYmTceDrxBphK4jilZh6s7eaoAlFEbRT9YRwLaqoO8ZU4xtWK789OQocCA4VBujVSa77cexoTb
xJTNo+cpTDNGN5ctRXCpBFW/4uKrEyrBvasaX0j/d7svCNnPvNm0els8TL11I6IZOMEL4iaGGAzq
wl3TAVnFk9bAueOK2KFY9vGUkE0pF5m1m+T5c/zCD9jZWjHn7CzfHCcUz6NAvfjCEQtD2yQQqCXz
1Sf1vRLGb8vqYpj6xY2+bLOQRtAOzcb9G3rurUAQmGlTh/QBSS4m8ZK5gvywdlrYmQkYH+WQ0rJO
bExzPdll5qcDIhTsZEJaXSJPRCkpiVfkCYLwnx0cevej/8ecQocfSZe8wAGWFS9SOzHxXaR8hIy1
+AWx50zuy4cWzinucmFc3fKsLlVcFYhN31Loa8iE8ZDl+8JJCnp/baG4Q4PDok05TDhYN9MDp5fW
/UOe4REhejmUX0s6LkZ1DSocro15qHUrpto93tkPtmA3DmQ4axI6n2T6r0XODmYnJDGOgqCxf95E
GdSTxAfwF/Yp+UnPT870PHgrreG0rILfrE1e6vpMD4NgocX1rEHXHBJRaKmp2Eesu01s5F818sDc
BfdGGDaDuLjLcZ01hAmovT1Zs9hLFgwa4DQ2sJe78jAkAn7G6y1rZLwEehK8WTVyPJlNS5SPK+Mq
9Onam2l7leNBjBEyTwpoQGafvdGRIUQFj/q3Ah6ZFj/Ht2vS8KHqtlekAms8jACi1Ow6GYTASqNQ
XS3b6cVQNm0nN+2aPACwlWFBf9rRYwiHntuyKpN3wCDvqjwdj8snYZEXiIwYXnjjtLtm1si0+Ccx
vPTMrRMqkBCY6XGz5g68R4smA81TiRoeumZhhEga/T/wKOThjHmn9hP0N+rFqp5Gsb2OX2V3W35Y
8CBkGKWQZuiikmRE3QPfA4YvLDcbuGNeXshaxKD97qLmUtvbYOSfU+GwIkPmTsJaREq/41mJTkWO
IxeTUqeYeF7IALxSAbGzFD8k8oHd5Yw1np7YrkX5lcCovmSFM3WFl9VhnkopEkrg7K4IdAUeOWaX
Chj5YY8DsB4bVTCujgjKniUWJusQrJZwmu4kp83rglyd6VcUrONAfRO1dzudpzEHUPVRCT8K7Nzv
GGkULx/3rgI9gAOaCWiH89M8u5Sp3GjFn8ReMYIcv8ABXmzRQm2jaBqAraxx6dH3kC0fTujlQB0A
Xavq0NYBj2j+xLLlI4QzWqD7+2kBk+XDLutoMYeoIdpBDg6xIQ097ZTkjJTsP3ftM2i1fhwBPFnf
dlk2OTamTWXPxabMvscXyH0LWiz+hu41U4R5vCEEN9rXaeL/8l5kgC5oTTKHYAnFR7u8jyLt/A1k
EPieAEcxJ9b3CXmPsvkNNzmy6Nut2ua4zF8fiaAldGx6WhZElyELXLpkiMClCrOMXai8aZ+vJAX2
5pt76cl7A3jPy3lBZnIjkG9tOZmtOZu39LMdVIiepqfDlwt/3AVazfQ8LwkruRZfBXK64/taPp/0
viNlga9gHwSLqMqNnE2VkgIz1MVfxLzoF16A5SaKrGKA8GrqjYFQd9IdnL2wuT/RkjUaIuGI4D2H
RWDOG1YOauQseCLCqhiLUJkpTKyQ/N3/FLfgsrfYujwd3W/TeZXPakhTCPy/E+CDGZx5B3hy5Xnt
QAGZ1FBbeV6TPJRiY2oGuJO11PjY+/ZhaSfRMqDTGRbHpYWQ1SH2a7UyouQfod/dgiQBh6xzrjw0
DIXf2k896tNdYqZQvMtafe83sGlkiR5Wfzarph0LgWeNXFXh3GkrLqPDhQMMOMOpYHpAYzvxvndE
5iPbyzd7H/ZKpJqeunnTSvVcE8+nepnrb/KwQKEQ2twP4KP0TMxjA0Sig9GV0mr+oPODecCec9oJ
GvSoahjjZGVMgL4fYAJH0GY7H9pjczKOppHUV+bO00U2FyvXpmfofqbkzlUahghVM/8fc35LVYGz
pkaqvzKLEN7F6gyumKx1zY3Zh/q2WoZ8P79SOE6DD9m5utM1jTBHaXkPsxMFO1iu+WQfS4DFWm5m
AfmAnt2OJ5k2viUbINKP6PE0wEpvcbop3+iQtouuSNC8OwCE276NQBYdDHXCv7mUIXqwsAOzDGB9
thklTWWkjQ1tlm18M8fAbmcI307/4QguddoQ/TejtYuYFG75Zrbut+lkGE5JrO5wMx1R5m3K56zB
JY8ouO+fXXyOLijI+GK3O/wimV3xvJzc1Rv9lH7S4K7OPRF2eo+UgnENJOLAoqBKdBP1g2TdtgPn
NtN6Rm6y/H0uqOB/DndXIlT2ghQ7XCiCe7G2m3ARmQqcoSQNZOCQtepRkm6fcOEMa/2mb1oykBI+
gFpaW0kGLOsOomw2sDXMTTDW0Xr0kxXQOx7zN7mAdCah5vXGWBqK2a6e57e8RA6/SUQ8Gc/kvZhk
PjohccQ2/4apBK/erGmws/C1hzVSrel6iT7CB07KKhVGd01F8zB8p4mGcTWo1kRCfRPmqyHZntjl
tI0fGDzyVxsj3VNdivdzJQ4OL9QeQdPtv/LKmNZ37mF794tfPC3vwt97rZ/MZ9a3doQfhHir7mOx
beOtukTKhJsvATAYF0oWp0ZkBFV1cEgRh1WJs+SxDtn9RHMOCX/jvsGcCGXhCztsV6o8kbSbt6iM
jnERHMzudexOsaDnAmnFU9EXpBXzulDMRNFA+cemSgtRe54uXRAtVf7NmQw1TjlPRSEpGZUc3i70
40mpa0mLxcAGYIespLuKCfJauWajw4Fgz+2w7EWCQuJk2jSa3yHJrtcBqJfXCfG7dPMMNUTMyVq1
x5QQvJdIz8uqE1Sm0pFs50KhEdUsEb8uLMbKoKa+AjHQUD4gLmMusNUB1fXj6Mnh5uSkmlMYOKl+
9lvphtOn5duUSRZU6x9zJXXYj80vaIqaqKPkhxjwCHsK5rb/KR5VpgZlzQ63YN0LALFbo2Fkii+q
/uR6Xfz/4z1QIwlJrUqjW86KtXFSK9Xhqi8GhqgeR2AG0CJnL1S+ojTf+nKXIcoyG4iAMk17T9Bt
jFhez0BmShg9jxavE8GtPzQCiemtu6Ie7rm/qxhO57bUrsAA/remUaP3vyqcHedVZMi1vT6TeYes
dyh7t/NeW+liRhCJ1ie60IrYGdrlXW/usmY5Td8mS0Bmi6/JqPsnVWWCTgPvHhZSkfVWNOT/5spb
jm0DvTMTgYfVvSjX4QifcUC+HqEX6v4+DlubRq0ctEg1ygw+phSHflqTp9NaDN+wnycp2JTcq52F
Zfycpa1VviM6hitm954ziN6yIcMqH+6/lJaCAe6mNrAZSFM0XKXRflLjVVa9+rFQwPQqpacSgyoR
/0umpfcQqdz8p6LDdjnnfv/xWnSeDSMEmO5mdsrwaEjjABPVdbtNZaT50JE+POq3wEV71umM9tie
uzt1Pn3ZsUZIXMgYV//+ErLD7Mc/iduKBm3pzliT7sXFsEU9hWAry4HgLkkR+Y33ReydkeRvfaQN
IRpUaNLW7LTiIuqn8vNneuYkMQTddQ9mSE+Y65kXG1hyko+c3cHuqWnhr1lvazfdxt+5JnNQhzz2
cwtAZrDJz/wHuJ2MNMPlaYEYUHNTkhsGVZ78tBLPAx/NEhq82P3EAX5lxdKLK8PwRZ+EL96xHLfd
xkUcrBctAmYiV/99MLqImb1jKgWlVaxg5EqxaIlBBGye5ZAw0xoOiSo5WNX5/AO3P6xjfkFXhdk6
+dxwFUE70kH/XlHewHqIiPEh/Gc1R1D8c8s9Sr/tu3UUh+ir0PP8acPvM+fh5cd+NKPmv5zKj4bB
qXiHNmAVBfBXrW75wavP7Ik/MJwt8J5agr6nvVL/2yuwqQ7WADx7ZZDbNhfYpRBpoipc+iNYh09f
GzYedoJuNOMZxWgnwcuTIwBgYgsUqJOAmdQg+ZsF1u0VSpuyb4xs9DXc2+SCNsqFzNe7MANvIsFA
7INOC11tdSQ2T3cV/P864y4YHzIvob+yzPLTetYMfPXbHPLChn0qcd64oBjDyrmUy79TfG/lNdwI
pLhIA7sSUEfNgb84GJquj795ZMYc76p6hynaqu6rNurDssz+FyP6DFdoxqXT3DgksJ9vV8SOTZ2j
ZfT2SClQ3xd79YuLCakC5/HOjCa67DF2nrRXaCJSAMcpE27Za8F7irgb3Kz+gSmsPkJsUNPegL2q
ShAUbMsdFwrDOjw1tqykjppnz+cIUHulu4CInowGEUWn9q4gz4sMlmZ8+ncIHLKw3fmCBtZbrap6
WcBCeZeaZdk4PbbexDcSofndzIcGGOf4dTuSX6VQwMGkHpfyNwi6u39HTI/YTQjWJ8P+bzKfBCYI
kGe323AOfu80Nqr8kgSjhDsxEu9W6x/HqVY+0G5XnlB+cAEdtnRs//Wo9zNHFK+X4uUKry9Az2Mo
KYxFx9ZTCy542lLsAS4fFAMlOSNK8JBSYJelRdebXQRMqBKxURHZ9ZI5ta95Hq78tC4miebNuW5F
rHDEYuf/q6PqECrsFfTdzXRzZ3QfaoNDqBLxG235JtM2joPKBVpHMcLgYczaL0ucHX7J7BgYjICn
CFWXY4H+QRh8hEf1clG0XKah50QBqI69xuxtPAp6qIivAUPYl6HFf36mFcEJ5M7q5lGCgNmS9CEu
wvlbwVaCaJdi2tcrVpq/exyNugX2NTporo0yTcJPa27fMSsJ8pxomHdVfpD82MoZ3oNupDaGoH+f
CHsGKzmhc2f/EutlSaNcpd6zQ5/yfHi8YscRV4OkiNhaWRjbOE4CohO9F5+RxO9Piujs09T6163d
BXBR8c5rdRsiw/74F5BZzpISq3FYhByccFnoLx2RCNHaigtiH3/PFyfuaX5DhlVSklIKnnzC7ZwR
IsUMiPnNFWYvcBgHDOTYUoByRulW92fVGo5G4Pz8CFNj27M+PTBHq3NQDStC6hnuOIUfh+4+G/Et
Zrg6psWLz50hBtcvaHfNHURvrijBShDUREbBnJumuLrs512F/OUbnz9ZbyimjtGqArceMcs+aprc
8Tz0YmrrBAHnSBdLX1B3hzQnD4iaoPPpMBC5sxu/RklAilF9gitKI/47vKhEk9htkCpsHts/MDZl
bEx1ycF9j2chKUkQmW7JJb47tfULMvGSj+aiiciz5Rn1gI2RP3ZEOcEwzB1U3fMqloorQ3zC2YHl
KeA17jzFHbd7Ylux05R6lFo2yisVfi5+81U77WRMbN+sBvkWH29H7+dIx3Oqyx+yYctQyP8QPuwj
WE3liDTgiVJlWBtWAIDbDSznwHxglcmjWHdpgFQ77SFlApz9jk7OJGRiG6kSoqU7PjDQyJEsQW//
TDVEAC9cKkI+G7IzecS3V+IJsB8b9NfJeOaEU+iijW4xlXPNieEv2NCE9aOjuR6S478zCVmaz0ea
Vk3VHXNdUVARrp46LK6E4gzaTHj/kM8JP6LAMIGLVgX+rkHvBQkweH91oiDrjec15acBNXCB/wlg
fA0no+190o1GbCPLOgTRVlhUGJ8zGlWIrNE5SdoJZs9XiBF7C62MlJQ1Nic5n18LQ3TqwpFZc9Fh
Pp7gbTMXBnYejhuY4Zyr32sGRt5Y/J5+pWMuTZRdcx9m4MZsdyOUsxLgAiOglCGOs0SFuNOjtcuu
A2rp3dCVkc/Uoorc4JqZz7EWRhj2Wm5C5SZHDO2dZzxO8UAOsptlVRKaTJLu3G2+wJg+tPOu9hdg
w5kFrHvC7KeJ5erycUhlp2/ZUF7nI5VK6h6NO97kVP6PQEeNNl2bJBDbMm65SjR7Z/aczD34SQ1r
5Jvh3PX52xvkzW5n4ZbO5mHVSIXfhxfbTfgyqXSSqBN2Iyyy9TNszqiQ8ETtpoo9f7vU7/79jL2w
H1/TYjM8eH3aa1td+IQVUViwXMG0Wo9meeekWkiLv2dTnlQsfMIZNkDQ1ujXC7dYHGGrkv2cqmSD
89+avc32j2C2gaNBsO7m6hCrrTDsGM/5YwlbfSpltsWuXYcuUIv4MdskRIYOTFkGP0aWvD6gyql7
fyVav2KbOfC4Lpf6yo05O1J4V7QCitxYiXwB3COWrGwrvs+s7U1i31T8TucRCCT46VZBldSGRJPU
2rTTNeYA9B9q3IwIty25MxQqxe8Pn1QtlfAzdMaDtOT0t/4bi7OjuUnGmLdDpN9XDrKEuNz2eELm
RF83b5FpA+Iab0BBRGx218HDh2FU58jAgMcZtlkkxt3E4rKnLN4Z8C0EbMv0EwYzi+TBtJMg/DWY
j6qI9QEiGuwcZD+vnJJajrZxRjeaFd8IdPPE34n0DKOlDiJExAa27ig1iDMugcmApUXRwOwLDMTp
01jk200xlJLXCabyjnOrTMVLkGS4QiEe3PHoplrxGfzz8YzXy7iku47I+p+9fLFgIhFLZfzew2Ap
6dLZroYVqnt2Km5vB6GSH1XdVV+7E2JJENrZ2R/X86YtfMs+I09ARP9gr3sf/bYwc1dl8AHI7ST1
JcqkxkvRfmyOCvFd4+VmlErLMNyCM3uSfS9nkDpfSa6UJX5NK62TEvZdrJVCuI6eCPrhwvNMXhhL
09xymhc7gmXCQuZqlq+/UDdT0mPc0h+xxhUhFsK6EZcmNkzYeEs7MdFakPSaVTNbUQNn9Bwl3PBl
7CCA6tu1rIQuVYRYwfgn9skD6srY5EOpG0yUE3GIUb0S4ay5LukfObz8T+tE6zXERoooZBFR+epQ
cqNw0Hbc7WguxARhlupbiVlI2JJcb8U+uC7NahhCEtvdr1AypBcbLyvPfyxKFXKbLT1Pj5dXZM4j
G0bgeT1k3li9QS4HMaKVGBCzPUTOZH/YfURkAKzabUBGCbyvAUdQNC0XGMBTIQHYiQvdFVMLr9Hp
ysj8qyxMUJDRLUSWzch2OQyguGBD/2AKVoCZn9ik648WU/uPVj6E3HlvlVKV4lSU+uUqmhDS6Pb4
fDW43+ePKRP+autcssUUN8GW71N8Xag1cHSKCWLSU+s0RZgx244tSFu8un9tOXceMehP/uoxCKf2
KQgBw7b2Aqwnm6YxYoai44kKWO4yZFjPKqdnxIoOjKCUybpEzDMmStiak0aNumvC4LjCe0TpL8JL
AEmelvCwrTDaxdCU8RLAgLlQEZKNKX/Y7adcbP5dp03+wv6eglTuWRb0gKuQTCNzo9hS08ugVnrS
XdMP4wxooV2R7yS5uIrUus0BEZDzMjBZnIeHsjQlB65Ztqv4xqMkKduAPlNu6MPzN/8Pxoz/c4g3
5nrSwdx0KbO/NN6BbwdBxvKo/d7/HG4N0il7Ev7UYIEYaom2ADZ8tkwG991DoSnc6MNtaF0Vy9/U
nWeVK5b7Q3SVZebglRUWz4UJ6z/FwBydKgYqq+s12dF3ZwtcArF/ZvleVIZnral7eHgF05LeX8xP
tce5IN1PVFJsoAh+Zcyoausi8Sgr6HIOmelDQgIZnToYrm5X2tfCmrZv1TY931s8x2t5lOwgVHM6
TpR+Toqlek2xRRwKMRXaAx9v/JCZAQn5f7bf+Zy+IAQck3ClLhEWMqjFXx18o1XAtgDQHDI78FwX
IKeiJaGa6F9BT/XOc4bwf2ZWMdEPttr0sa9PMMvTCinEoMVAIx0v9PbSETHUiCGeLNZEdOFg7UWR
O3iG+d8Pr+pISGbz6bljg4T3B/lPpp2luVQRKqBEHPuWr2c69YHK+VqsnP9myFZ70MxhE5tYY/1b
OFw09biTY0qqyDz6FJi9MnZkzx3HB1tTfGRdJM2UjIOBsv7349hi0L+ZAjSs+8fctVXuHQhwZRc9
sdkZ0X4Sqwi8EoxHDyGhDVKyabEIE/wbSGAcIBILy+1yr3j2DSE5OAFvbiXBP7VfHfzt5+urJxtt
v1TjfpZ7/aL4GEjDXJChdEuNh2PIYLFxn1Z3k0oWvXrKFPKprTGogsDFp/66qWE+F3XkgXwzG0ML
Y9iN+9uRZZtd4W2mxrsHl5gLeIXp+ukLxO+ZSrydenqQlkdRPPBM+DugxDR06E5vxmihHhcO2QEN
QiEMFXn3zL32tXJpZYHmOIMk2ujiJzwfaP6ERUVEyYiDFxbjU5zom+b75iB4jtUQ8ThwPvPslaUZ
a4DcJJFK8SZKQW0TMI0HLTyN4G+ZeS2kej+Pq92eJAcepjCA5G9fdz90KtCRIibEnLz9Kz6+Jdfb
fROX3UZIen9P9doMkRsB+L+qbAl7bnsFcOaKe+y1Tq/NFjmZD/cLoyWfH44matRPBSZ+O21oB4tc
b6Dr4e9nzhCud47jMm69Z5D0+7//sZtPjV5zBsIKpIDgYg85bIHl7IJx5SG68dpvOwJr/VF3dNHN
VlRos7jVGVNycCHm5rKQdGs+5a0V5SE/gUA43X03WTk/HM6WRzdsovpnd5wRi4r/64SpjFwtgXAW
QIW+AKV5uocSwZJBMIBL+gQ0yO51M4U8e6AyVPSY9tpdt96iN7rR9p6e9aWw/uZgt3wJAOELex8N
75+ukBI75J6zDsblzab1KraQLusUs8VULM5JOMO+mJMzLR7iluBwJqDtUR+vAgK532iWCdvhNmy1
qEOHmJ75/sYdjMH8Pi7OUDIogXcNNZ7yDeN6bUpXZyMTIbehd57p0/OSaT8W3j3bs/OjoMDcQLTv
tylFvkQhnQp5CkX9AQqDia1SP1Mki7p08sa1cQOdP35QUJQK3nnWxw/oHi/+YmM8uNRPdImxfnfd
vczo0q0RRSnE/T4gIMM+qMpKU5fEOWq27MOz7+vQdkLlC94arD+brH+woCB6kjFa8EkN0E1bxnjm
4oHk7QXOuQvyoMc2aSQuMlUIuZOh3dxCrCXitOxtCll2CD6t/A+xm1k4IV6RoDxwTjo6NR9wDYH+
p+cuVsGNtyenBunU3HzHYzk6/Wl5jVcFAanHcAVImVLP/InWRSfyyG28W/IjThp+TSg4EN7HIHMP
5kRmxfvXGsKi0WcgOibAtDDNuDABKxSw/PrBuAx2oOwvl20Kz66ZShcyb5t3a7gPDjJkvm48Odcj
n0YHanQHC+ME5DDRC05K59GXzcPLsmknGaBaimHLXyEtcq/LQj/Qm2kygEQvaqZcy7OfBCcaQJoj
48TpAlgfWGxX3x+dQe7MjmkI0gtAXS1tn8tSIC555rzKmhZKjMpj7nYZkfm4x++X0HorSGQ9IvuK
zV/vvtgDfUCCN1noJ8Y6YlnsBxc9HVG2IF1/7exW/PqEC7AH47c45hlvUFdBYqaCR05RDyzbnLnx
yvcndYOoXkbwqoVrpBZTuUjChRvqqXhnjJeWEhRETV4bgqJsO0GvB9CJfl/VS85e5R+YkbsuNM5X
QhBKpcjfNGjJj1Kldw8L4Hvv4C11gXTff5yXR+7LQZ+Yb7sVBldBzjV0zRRdGlC4+brWgSo+SVsK
73mQnDggMwHI5sj0RhkwsyOb/J3+vLcEELL7+f60wSWf8U4VgRQMfHW+9Qp5fNX8rUP2ASPENU3V
IlQTWozVmamedXSv5Q3e01yXv2KRKUoTb+oko2kVXfANYVHfirMLU59DHldg6Tx1Nr1dCqRF/mk4
8yYehFGL2rkvKAAMSyu/vMc+juOtd7bWM/uMhYyNZoMgYSKMUPGb6zy3Z2d3xmBfdEx+rHGCTlQZ
29jwJqCmdW+mvnQRD80cg11zq1Favy/BpGArlBGOMzoD8ULaJ4xCI+HZP4hBNSXSfVcKe35KSyHb
mn2yjzWnGHogf+7kikZnwlwqJx8d8ftTlGxIb2ECFQaETFz2zoFvkUZ4ES8yxaBn9GR4CzwPwLWy
8YlslcmJwyX6bUNpU9i/ZHPEx/xqYT9MsguTXM992jidyrlW+8VbElJQQ31Kzf5dXNHoJgKgjAY/
pBmnsLMA576TTSkYsDdvG4Hq2taCtEQeBTnSRCLEg5zicu8cIB4y26AzT6Tce/kube4nBesCG54H
wx23xjKht3g70OObMEZEk0xwznXHPh+6YPaiclxh98Nj2AdTgINkiDLJ2QRvGjuWTnmCn8sxaREi
pwsOpCfZ8vhNLg68kPLVn4Wr7fU2OdRoj3Qrm/RXBwX62S1+ZkexWV4i3NfmzgREENDRfTWlD3nu
mMXZ292fafICgjOe5fo8dZ6jMmY1t/gnr0SYjPkEbDdaw6uPIkHhMyktRGKgWOtJX1V6+lF85B0i
6H/5Cbp6HP9lXngkik/O5c8XGUKbtWz1Et4ad2V2rbmeGvP1rYyKG2ydVzG7EMj6e5jn6M99coft
CeY/y+16ppz2DRrnjSlgQSKwLgbR7WEfuV4UqVe+5XwzEr1aIQnD0Sj2Ur1v5ZCvt1Jlbs86bqav
rr/Hufq3/S8vcmapGB/0oNn9t4AhyRn92/rV/9qc+gR14ronFnFMtkRPIUo/ipKJoNHkUi5kVnVS
EpAtYhIw+oHZ73JarfF5awZS/ESM49hU6OwBOdtXiAkzg8n6juSE1gdjYKNhMJLtUj9si5Qy6v/D
pKES61AhoFRyLQElo9/XE7K9xZajuVy406rdpaGD5CoK8iPB5bHfrc8f8cURuAMfDqpEuruCzUvK
p6+A2paAW9KIicTbClofF+7tqDhtC/b3Xg2ZYbCsdI8D+UB2XewxBb6LQ90D77kjOTRbfHiOnm86
6TGkJd+OvscYPxSwbxvAeBhRFD92YV2pfzEUeOjt480yNtGmB1bgV4FXmGkg561yP28YlwRhuASA
G49yqVRfsHBxXPxVyZOVXWs2mNXmvo2cWjBejy1llsnoK3jBQK9YgcYtDeBMTW0BmxhMXLV4Ze5p
p9zGQ3ug2zuCd1L2PSO2Mpzuq4kFUF0c/u1O4wC1XAkLq4VPr/2ENM3kfm7XRLPAIU184HJptrO4
f7fGIEWK7Py2i6qrWbH1u/ttoHuesogIWC+KFhqrljrOaklSJAotbJo1a2dhdMTJz8FQ1M077U8y
JKxIXO2V7Z+lC7ZqTWqdSlLuHxqClStyhQlUk6z3JqCv9HYXmjMlQjrKlhScLTDV1eORVJVGmcEj
tr5bQzMurXR2f1/ZHB1iRm+gssQ9XEajahgsDj2LAqNXqm7C79iQlBmTa5rNecOn1O5Ifte6tsF8
thpqQVKA1ZnXTIBcS7R9+hoTSOWYQYEGvYsELDa+mry3fqWTUVTCL4U4UjABSFb+E9448PqMnYw6
6vtL68cgcn6OJkyDfC3AiRq97mKkymrE7VxEkSxZgWYUys2saykcxC9h/vXhT3QoAdDMXk94fT7G
m7DSXCejNaC+ONzM9VyUAIOwKPGEbhMBGHAsNYMbiYF5CPZmi9szqh/D80yawVnP7veTDRWebuh2
nd4HXGtiBZBayhSXHkPq5qOFzILaWasAf7JzATZUUYpz6WQrE6GKX3OQckEuIfNg2Y2htoQzWs2H
lgJl1+nuj/20CoHFYckWsubRj7wQ2Au688E4n3xfUwGMFC/Tq+EQlQi3BOP2SXf+ciykWhYIHUrE
wo9bROX0kzjprCCkwvqWllZ/9k+QWVgO8xUJ4x6ZhK5xodoR2jl+76uDxVQnNUn91Tig3Hi4ZM5p
NIx+VAdZc8D5c3yk62TCGKfXv5Ndi2K2ZGn5Pxv2iSNe7Jd6/CXtXC8aW+S7zZUMrgg3BZcHsyf4
3LPXkiCeBvOFmrxR1R/MMu3iSTAV+EYv/OmNj5BtpAjlHqJpXGtw7AN9Okfbru5PaOXEIx4JpB8s
34+ytfLLo44nzBhHWCI4MYm42LaTxZUcUIApFKU2sdSok8CpS6/LXeV6UZMvR5sZDtjHdJo9oopN
6yivuIUTDbN8pfJoecgh/6ENZ7VHs1qGirs+Vga1hzFdMi0Kpp1Cpj55mBKwQ/+TqXUyegr1a03F
YFrnu8uUcfjkN+OL+twLF1nJPWi1CDMNiEFmPyxWzlFAvApvUqoBvhrTZuIH79mkBiHZ42LJRm9Q
Jihb53+gJybp0BBSKpitYIw/+yNTTWJnm9PpR8hgeKZ/SaNsL640G/EaFq4WPuwnz8jy/kjlKRML
lZhKNYWP4oPPAn3t8AlBH0xMCRHdCRBuMWTJcvA66lSD+Zdc9XXZBHJ/Wr8xcFt6b5qPbAMOONsx
i3KeeztKBui69YHT0KzNI4AWrLpFb+ZUlAJn3VyVbjt8sknBFSpZWSJEnVYBIW2oA87gPbV/IyHe
9sP4HD1ErnCJF0dY7VoWlC3Cox2ejZx+NWxRwjygbAA+fAi9p+5rlbr1W0ET+pNPuJVTJwtk+dMB
stSpQjZNATTmBpgw1vMGn5oQOmUa75QQcQX2V+c2WeCz0pDcwKYL9Skhm7aGw1Fp2oL6iHfA7qOR
T+Xwr0+HI/iv3cUDilmUI93o7arYihs2vc404KqwzMHE+rNBoUzhS9GuEuSPvIxYYtnARbWWAwVW
A/mEtyxpscHj0mu6pm6EWjj4winN5rARWjdOWG/O9klfE5G+wj0EJhmU3zFvqXWDATRO06jAXAX2
sI+Rl6xTEcQNscnQTMo0ZdecbP6kX7RAK+FV7JY9uQWiokhS9BStMYZ6UdfbrUghDShoJ67I/4vt
KqLY4w3JRjwQU2TCA1+OdipP1HUqYqlyruA/Rtb5CiR80rQ7iv/RSuC7gAfRAYRYS77rnau6tCJw
oFSmfqfdsBKrJRD/K9NTEM6KlOHP6t1x3Xp1bl++qhjNC3pBJXTk3zKWcIEGyA7LjBfNj76x1Wtm
+5eTIbug27eFbnojg5QpXB7d05hyXQp8d6b+1AVwqKUyPd8TxEGGfrPotqQiSALuOxauc9Ybe6AL
1xhLOpNSY7VuL3TUgbB8Xfz9Xf4kfvmApitfh/mRqJXLv3X89Uz+3yMDOuE7JXXyM610pR8PKx8f
ANzn28UW6i+LxDD9Cr4pD+Ry4SAOSbIF3JF4Xwm85Z/4TIPzF3IFbIdrYUe/vTCZTmjN5jvVJ0RS
6TAQ7t8wAAUjYHgFQSXRZQL65EcAca+gC7CCfii3Cfa8WM62WgSxx/Fnw/ZOqa/ZN87tF23VqWkh
r7bkgnllDvnmX0YV3tYQmozCi3DuC6LPVeDZ+XDdJ41qcKFB3OZLDPLPyK1rN9dcFsPdUMnXiCA1
h3xLAQzi0rUtfpjzsMmWvr4t1YtRLIanRdRJSWi9zP1eTk3PNQSOKCg+Xw8SPObKIDt6XJFFeRNH
B2GBFS7JUkBuY7s6x62Xxtw8/DbvJWjkkl83UROPCxfo+3K6QTzOFTUJog8rtjx8A+aQiH/U84KP
G14A8qCy+disQRPsR7eYpZia8jOsUo1nxKzmJ9hHNuHjhqEW23su2qfKcRdC6+6RYT7jqc2Ih0ww
2Ko4sa825Ngb/YvVhQHiYgxuOqK2P9yryj4CnQYG8U0SXXBGt7ose2XhnkLrKLcEBCmLOUZXpECu
lhzVhLwYkHjakdgHNAOrLZcqqKO85gOAo8xR3eoJXN/zYWi94AgxCPnLhhHIA+dwAXYznX2nZ5/x
6nzgLE4bgtN2ntcq/lXOm7muTJrzOZNrFOHQNSPwB+09Y/IVrRo3wHz4L1tQGUFvhv4U9I0L9ZsL
gvoXEfVie6BRwhGzyDGqgSNTDo/Ydh9pxM0ZsXQhqpsZsD2qr5FskmiamB0/8h2R4cFNjjAlXzO1
k3u/uixHNt/l3ajnQPwNi/BwKqUfJKBjsh+331SlcWY0nb3oYV7NS4GAZ9JvrlSBCct4oiYnKKV9
2zO59l+tTdGCSi/Fx6OeaQMSxqzaRHe0tvGTU2LhkPBwGWRikFbCTqjBD0ptwpaCjNe71gUllNXt
kB26Lcow2Q4zN3RpaYu8flBOiQ/SSvph7e1At1GA2xP3rvk0yiumiA4DMSSi9IWOgz289Vi1IHu+
KjKOTYdwK7TNzpsVB3jVovg5ZvXhFJOn0nYNmCfjd8Z8gG8/MDeRk+2kLZbsBzox3SQqKmpQYL9u
VtCmQ80/EUm4F7r28GqlL/o8Z30JAnyTiFZFTVdqpPjyQuA1k8Uaw0r+P+p+QxhCYyWUzcaItMGs
Ijdakb1he+78ztGB9tof55X5aOywfggnT/e5gs90GmtOeUT/H+XeaI5N0RnnYhxOH8lqfwP6EG/S
i3IZ5tcbiljs/hqLvJAdkrfTnAwHr4UB+8qMb/K7NqZVceAwJvwcVEdrW64eYUNlH/hMH2Bxzzpz
wnGmc20DvKUaEDYxmJdADY+7juIb23t+O1vochTZx0LPJsX1zHTZy+M9dnwFmTExfMcijnsrsOX2
wOJfyRudtz9/lAuFJIAcfHu6tbRu+G2y/NorAOaJUSf0lY8FSHwmB7MYknhLu+QYT2BsAsQUx5r8
cGDpQzvzsOEc45YJ1bVLuFjeKf8RmM0BALo2R7xfAKyeFXgwK7ywYxeKyuzUFhP79O7+ThySQKqQ
41w9NTYeV6h/wbAekOuQ908Fg3svv74d7IXa1XzLkZLkKdjwjry2gYSA85tWXNRwoVqlBGgsqqiS
9HBPCVFQDBsYuzqXnbikc0pyfkVflnat1qFSUQI3mvvmWBGTxWzBJzYUS16FS/H8jgE42NGgTISL
efFx68vMi0kWA6+qPsrLwjakJEtKo82ulYa0qI+MJrAC8o1qRyzMo+pu9jV7OuNum4YAJ7w+YDzC
Cyss3b0lFaBVW87LuURuaUa6NGK24uh2LGXSRxAzJJVhIyu4e21YGBQM7zKWOM3KJSIMzctqjtRT
EW8B3gtfXt+O8ni4VoO20+Mfw/ppxGPIye2kTS9sXZSVYE4rzx2HzdRJ1BW05O45/u0BgVNVYF3n
3AIfkkZHB4aqaQ4jQjU3YJT7exPqnWrhhhrPBBuxdSIDncIpytNsYaAT2LCp9dOaD72Uuz8kl4gJ
3y5wMjR5fRc0w3ybNxotzwz5tacTacY3w/AbOYWlkiOsYyAhnN0QsXMnumFIJ7kS+ueILYhxHNqJ
oUsV0MZvuqdmhwX/3ULZbpaf9/izUgrCHrnUUiYdFl6ra12dBfPnYX2xzohl67HieT7wKFekvECI
ELvzEdmUWSBF3xvxlzpgBHY3aYuGh4+tE2oP2HToYkQysq02KYcmNnszgVZOvBYP26EHvj7gMgd6
FNPESw1BtQ2oHNgpHL1uqJcfOYfppSU3dm8ZIlFmSR1AtaF/zQRQITMza1OISg3+nf4eVkroPAnI
uCsAbh2mLM61FpMqTsXDfuX5nMc5tXqq0mgCAjFdSq8uMa35PBuBrJg2lltOy7GzE5VvMwt/FBux
U7sqp4/VwunrKiGdkHJcrhAcOagg1PJuo8Ty8AUY7xCabW7GZlO1HqNfwkQMkXoqs/EWFVe4Z9uc
sNLFRTug6xKkwEvvWxT7OXYMulvgu47mt9HjVdpWZeWTgWX4IyCJDDgmYzZTI443blvKXBlqjmjI
RGl7QVNsMOSTw5yLDcTGfY4w49MJrbNIpIxfH5syweT1yavMmO9xo0ysvdk5xC5UfNRhiILBbj7d
s8Xl0hjcELQy+LG6+bT79Afn64wCLBiDyn7b8fU/sRaSpPIc5eeNB4o9IAoxbIBTc0JrDhUU7Ye7
UQ5tIs9FgsmrqJfc564eullVtrRdrnFrG/WYWaYDLWU3vHTZt85Td0QwHWS6nmOPuN1Gp7cM1aUf
DZErJ+KMiBSiJ9vVIaccu/sLDSYMJAB/kShfrWFhRrdfslAx8JnF66GzyhtapP4IU8qTsYJIk5Ug
bztu7zpIJfXmUmtgGXrUcGDzFjM94Dss5bBZA9RLi0UgzgsiS3cpdy+zLepAVM+WouC/36XbT1o7
S8c+tqlfWtP6udgwwIajo3UCehmB6AvpSUJcazf6SIM4xCq/Wmy8F9/ZYnMsj+BoZW6Wl+SDd0Z0
49DOjWmypdCkV9OYrJhsgr3shLU+YSPYH2h+UNeaqoRxZnL3bXai/fimuB2RM+u0KH5G/1FYnFng
sAF7bfj3bLX3q2op1uFPaGoi1qG+jlhsbOKs+lMebFvaQlgNtb6t1p/arF21CkcHqtBPCLhuW4Dg
5cOuDD+f3qWJ+i6y4No9L5/1uOA6Z2OtmsnfIcPTYHPW/TCSJGXfPHnNY0xbUyj73VT+COshI172
OSdCm0VdwsHz8dIGoHesjIYRQvrKBEdDwFC88mxrdH5HOWTFz/Hvy0mC9M4rqILDqGYEZQG5YFNM
2HelQsdS53WpI6rN4Gbc8ODvLMrVW/TR/k1XyLK/eiYqmvKof5KtKij3TzzNlfAAhBg5jE6ZXVZA
rYEGGFGKxPuZ5y+Q9tQOa0y4joaNSeiL9BXwnjaWUMY18tXqSoErQmUCTSG5/QZMvV6RF3sGDjo7
K9Lk3PBJHohtnTDwI0WKtWO3rGDEe3Vp4fJRJ5h9rvMywR9w89xIdlbMeTEGh6cX3PCzF6VAr3YQ
56NRAfglDxuprsBqBsHvCx4W1l3vZYjzhmo2tzsZFl4JnnyhxYfDSAFt5K0iAc16Sh/cw8b3kYlI
roo/qM02lM2S/+mwcJgAppaqUN7xmaGMeb9wT6lAdpasY3N79pGqLOaROBShxx0WoYOkz/zRDqg0
tqKTzrnVD5QxxJZx2gGZ89nq/ffExKJ2FZ6JhRdIKx8MBpodMDs6SWPgzg91ozL7YuJzVZWYep7U
SM1RdCUKPnQplUC2/7XGKYVj1lvopwvN+Z9i5OYdAPokIwP06kDQLWvOKuruBLRJxlqAaJ8YUzeH
hseM9zwbu4rLJqZ5enkiMGhqN8NFZnEWk0lAy6d9ilzGiV91rZEbj6Ds8n3LYQcQ4G8sRR4qk877
7gddxLRxA0B6YnknB3668GuuBV/ggfX0HbZi9XdZvEBQxT8iAdKipd+pCb7vWrv3HqEALm1PgKcx
GnoIKeKzJM2nzz6FA72xEZxJzfbgbovZV2sGmvjvW++wsW88UpBCoor60Y8LN0zwux+TVTVaUqll
4mkJ44KnqM7ibuNiB2ZSZdVGKvkKidvZ86VUdJXJH8XF3Y11r/7Ht2+ATFzchwl+3GXJJ4b/B3sb
oYIZ3xYqj3loKObeTEnBHaYnguBJ0jaPYdnoGWbcmY1ERb8nnYjV+fIwBikVMoClHBEA5ZFigeZP
V70sWKGLNSgrc8XvS2YK6yeKnR0jBDytRvXJNXTr7mSak2FgjH3QeWGwCya0Otuub3Q+cZn+5nqv
gT9on0+3CgJJ8TylP6i6/XQvH1fQiqyM2g3yhA/ypVBbWZLfFVfRPxhwEgz0PAM1dG2/yeLV2wKU
dU7RCgsVDdG+EXeMh1mS1r4TZXKak1MHtAZWeg3KwOqhVypNl+I2+XgBgvU3N88/ignONzOFTD9v
agPCrCMlNkYpQA30Dri+gRPZL4s3rUGKYP/Eo8kZ6IN6iPYnMZIvV+bcfWuRfmHN4jXeovsv65nq
iO1LcU4cLJomHCnmq5T605MApMJPDs0ClKFCmsaJ7DZZdPkk7C1e8o+H9GfFCOmh7ZbS8JbWEiiQ
50bYMbUbbKh6uawiccmT8paBL8RIfPj6v4NRbtLUB49k7xQMQE9bQjrnEFvrHWLMTyCcMRV3A3vl
451ZdJO1zaxWgPya0Nv7ak0cc98gVPhNjevNx0ZI9Nr6nuhazKZlDBiVMbw1c9SWFj+ZYj5FTWaR
ajR/gjelOsQIVefDZN4M6q7rus25ILOd8fe4krjqEOI3g0a+7aivx8JZHkh3a4zKfHS78UgdU9vf
3KNSK2VSA2IiouuspVX5J6pwZX9iJG6aQGcsQX1E7bahYEB1zCLEfSF7a2ShUepGLNdZ4kLZpnXa
dEJFeOAANKQBMKqMhQRAdZX386QO4HAN0L8YyDgHsvUe4XvP9Fp0lQPYnU4bFTYOYxOO8zCI46hp
qVdG6175m/Y4W+qjbKVMour817ZvGkWMOce/jaHHWTMWU9FaxdpSMFKa3r6Aydfd/bSRu2lU+xYK
jT/11etsRR+ywl+DGupxA0ucfu50szfrdfNHmsAro5d4r57OR74IGewJJFaNypueudK1NFfPvDdK
r4+RKjarf+R4NwJw5RWJUNPiHaqSD00G5DHRBhChBjspOwKJK1RaheYWtczC2/McP6jEdmP7aoKq
PpWxLc0YsE6hyJZ8i1ZUS3SGX4x1Wt2qs0eJLJAqA4hgxtDPj0j8sg+AYcKA0rA2fZZsA0C5ivbz
MNt2wFnNNjwnXlPL2dymzj6mZHefqucawF3b+ho3W2wH4q7y/TaMgCqjmdbtNEsyQkONI/3wPoV8
hMYEfSudoDkxCkGuMuW/SPs1SWlhhiTPb1jfrhazrroO43XjtXdq6PUjlZln1AU4hWSAdAhZp8/B
j5u9YhFh/2K0qhn77s5P0SmS0teBm2uWU7xMZxlEwEtMM9FjBpYTDfxA2PnTq7LS/2+q12ATVV79
9br+ixxS06CG4qZezqJ86xXjRq74hqtnW/RbFLR1mRIgtGqlKFlrq13qg8DUzKmQo8/3A46eYdDi
G+c/tAQOEnDLYFLspZy9oYp9iKQDz9VXdzJEcnb1wxc8GaaMMZn4+Wl/7p01HeEY2OVdpGUiGgAB
xqMlbFyxMiDkMLwDfsOKNrrCvrHrBf8vysuJIGm67gWFqWXozvqeqgMAAwxkyJytct7JugLT/xZC
44kUwsL3vYE1GLF/tIZdPktARaLZpnud+iI6aL6RFPo+Q8ms9g0lkskrzjk0POcXx+d4PuGOCp6r
adpl8mgtk+h8R4w2jpR8aoUAOl+rFZbBW87Vf/0Phg5szcc3+I9NgF3kIJ4zvFHOTVa5c4NWfcfW
V+Bub/OghXUCDFN8E3Mt4CXT3BPDLimJAIvz3vK7+Y1sWBsaXZd87fCes+DcRzh01l1yWz02HqL7
RpxVx+7tQ66Kvc9zQnbN1ZUy8QfFnY5eQ/d5T9C7zz0pY6N3ehim0qxn2X9HX1LWPl+S+UWXCTic
p/zIFqjMaDGkNyDsgwXSZDSwhQzxIbwcmbE0IX7Is6mfdINEEmgsf5HGfhK5Ij1pzQqsLudtA5zZ
rch4YowgpVm5+z80k3b8vs6qATuk5UViIkUR+pBftWqxThxUmW3/vQn56YEfSYJmS6SdgMG8ErwE
ajIi9kx/nBFeYp4xhPjzGuXEr2N5DJmJgS/OXZUMQN1vVe2jsxFivMis4/UuUBOijcQkjNdU+hqo
39gFHzSNoJXnzL48bkHhu6CNoV2kmml2tk6Tp71yzOXxpJgtjeco3NM/A0xZ7RJQ2qEOc2s7ckP8
KhzHU4dyAMLUo9FH7LTyCwcT9Xym9hEXire32hhwemU75tshd1Uw+1CHqeO2rf/PfLNjIqY05DH1
97P2XnP4psmqchyjlB/dJ2lqNzvhg3onUfsZUmpCTyqlyWErxQouzEodZnD/+Gcehp93YySMCv/p
S06Egg/qGwd0lfTmxiJ9N0AMaZDk2clepFwY6p8jw5TG0XduHMBKsFxMDEweinzi4JtSPptfJzUk
idKgvL0myZnBP4EuFNV01EnzaqY4fv0W7nX1Zslr+qnA/hEGbEMgsnNxOwhahk6poV9wCK1O53Hx
2xvrXiZmeJQfborl0Q7KuoWvfmR6meQiUlS4aNsG4TK70aHiVvSQJPKMY80JwTZ/wKFE60s5vVBv
jzej622Z2AjSknkTT3RPhzX2oH1khE92wPwOMi9bS1SljzNT6fjVQSCcRE8UHq2FjUKjQ16C4dCJ
aU+p7IOl1qjypqvyOm6n+q5p+EWjPzDJuEF58OfTkWvWbzheVEdI5LcGBIKDycIxGfihu3hofJyP
la8Yyf/Ks5MB7fMp2DbL8DEoebTLT4QnZzCo89uMgCEsBH0f0R8n0QxTeaURVYYsQw6nOQvb5tQ2
oaT8bCelzamH53/hF9/Emd8gMFgcQiER5Mi2BAdA6y55ZmfdRFamGxAV0PvQQiROO2NbS1rpgpWy
z68Yo9kZgamVyfSFY0AQwfPT5nS7Ny5E1zaWznROS7We2zLhY+pFTgFIaVWVeeDQmPxIr5XjNuOE
jDjy/hQlMgDvX5Og8EiaGHRBJcahQM09zwV7ZjVgC2XfFhOdHtWALjAItxf8incsgHLuO83hLOIK
oDmCdVqNXfalNIO3jmdXW1iSIANFi85OMyEQaa0eREPilD7BolEbzhQDW6CJQtb7m2+9THLLeCBH
wpJfjEIUCqcO861+UIvGwe5gALmK582g/H2uUS9uIa/2+xGxmEGC/DjWGk6QZ968Gpce+EIcjQKF
gOS54KLY+v7FZiMKquINvNwteAsH6Mgm1+HNfFv+I1PP+PUu5J7Oe3RhX5DtG6YdR/hk0jf6nBhu
sqN7g+FpihV0Qs5ILQW6/IiFVGS2L7QT3ggy9j8MEmbdrC54KWRH0GWKFePwvuhQw9Yq255SFq3j
wW2pkJGDJ8icY2gY6aTce53VFSI7UDZYaIGv8wUdtzuR82mfCGQ4hRUKSmS16OUf3sZ0YRT8TZgv
9wI+Vrfa8sjZ2hoK1L3zT5s00KkI1wRVySRen0cSXDrcyTR1QD4aqXey1kOILxUp74tcFr3RC3xG
8aM/KNeXaU2inlwZbVNIeY1CUw+XXBmGaKFMqGadcAXKD7RC7Rd/PiLv5CaR8LBXveoBN8nSypUN
i6Nou1lrSm1sZA/KfmFYt1fk0r8ZGkBSIXQIzTuNPU2b3YwSmu1etGDWuLrKXfjOykdNnJqGFYyc
QRx4UZzjIpfW6SHqFOaeG3RdU3I2jaBQbnOozD2ATmtrLPqp3WkX+5XbxluB2DfhhuMJHBZXqjdK
hk3WD3vw3Np/VQPWntYvgNVOKZOu94La+NlDdpZ+h5pHTY+czr5CYAWCMo0Pn2qPo3YQlb/ziPzY
l3ADZcX5ZridLhR6dl7NWTD22gXxFFAT8aKDf0KXLtaVcZwr2SX1j3sffepa8QG2dr3EwR9Jp4iG
VyE46Ax3ItvkGFWBEce/MUk5bETaUvaOQG9p66x6/2XfzgLx8GvFHapbiocM/yjc07nfEtg8X41x
fVi6jT0pIWF0cEXC7+DyDprxNukhS7Rtj9GONNZ2GpLCbQCo782orvIrnEcFiNi0ZmVHp69DXU0i
b4wb0ENTrEUnHnBQOKpEaH9+QJpnnOd4jAwLr7Rf8rPLVG2C1FneienONMKLL/WPfKJvA/w2bm+2
dyZFNCcvtCK6ASgSsuybKPL6/KOtLmEBoCxkeYXsImmIsldpINcfKtXm0ryX7fK6XErZ/Qnz/TRj
X+7YmlfxHDHYk3/urVSc0KX3fSzvIPzD3qVyffo+z/Q3R9F2tc9lQ+je/jdgQ2A/ie6xFVxagcWP
8SLAwYg+Iq7RrDdQDV+s/mTdDDXt0DKO93jN1h4QVxFCYfG1OoEHZ4fqbVillO+9mPn0iZppGGSg
JIWRFHOX1ru8FzFx1t8K9WqH58n/vXsUOICi8GRDXyExRk1Lzwtk3P2roTwDbJpv+ylPhQdXLlra
/W/xJ1v5q9jxg3v5L4qJdnxoxfSN8WfIGJzYIzQDNoJ+NmA1pD/138HdjKrx3zg7nRyzBLhFf+T9
UPIqyWKE4E6Z7+ZWcqEO6zCPKh0v8ipKUDwUviJUijiJZlZAaRZQWkr8GkBwCUXk+3gEvjvaClUi
sAGUrzbRt7iL48GBoc4UKbxxrrhUQiyVPAmZouIDh1Ij76Vn795SvJr95ZstHfr5JYN4+LZtPaoI
XgUrGVqpxOPPpNDiPwbTX3I5gqSqsZNNEZkVJsTwagig/BFZNxkRib0HrlRpn7SAM9e+kOqSJTm3
5H87/AGwePyJb9wpVedWv+j340XfTfLfxQPvkGR3EjSiac1fZy5B20iI23Dw5aNrAoeW0Njq4Qfk
wqAUVeG7147GGtMY5HfXeP6wMMOHQG/i4pxD7/fYTCsI7WtJnXhOX1nPUd3Z6MXEmUGHXwCZI698
OjbwIEgP1J6LSbcgaE8E7i/nNZ+1ztYY4zkJ+lncSHOq6w2ZdNN7Y+91SEkphLmmVvtBTuvMeCcr
cnY8sm2PG1evr3TTw0aSiBFjgZCHeOuoKCRq9G7736pnQ2KinOGrM0RBeNDvf0sFxnWiDnzYonP/
tUA5GjgkIJLDvuMDNbQh2+GcEsfJfMI/aIwv+BZvJPCzsfFXLX5FGrXuyQrwuaJcw7kmUo/fPam/
aImgCYREtwEPJVbkTiz1ohOyJn+4LoSYtaZDvrahpJkWQkGuiblWeBpLoiv28XbJkCPwcegrxrAK
3FnhJjA8brNGZ2PP6ZfKVR3feDRpNpepG8Ib3K9MKsDJMihiIkJhBfv8zkQoGe7XvGZlFDo3BQj2
MnRiSjBDH4BrPY21iwCDdcYMiA9/XCiiOkSa9iNquWwSOCBSaZVaCRcQ4NJZU1qMpU1FHgOAxidb
vMQKGftjKArxvJgwDokPCfSR7lXkZvEPtVJAgNjOJO9G+X1rH8u4XxPVstFHeRYw3kHJ1RpJtQRF
fFrrgQk1kCqcIPgdm2iGCH15A7zR4Ew2tMVQvUMRgw3HN/x1RLfJ1v4cgFUwHzGQWhR4o32wxp6v
8p+lK978uRB+XIIzR74BNDtw8oDBjsvJ4ZIbkDgN03by6XxQ3fOuaq338FCoVPvsj3cLUw7mJ5in
nFvWGj49ZW45EttCeYKE0U4qqOT6fKJPOjEHCk7JG27QrUnexJuAMmAYqTmpZ5G4HH4PazP9V0EB
h5R9xqEWNiZg1TSshNdk978Cb4KWkxprXyDHl7uV6haF2hIDSMu3EvN4RZcJEDFkIpgHX/pSNWAY
CLrGIheQQkpg16j0q4OsnsAE0a6lcubXHkHQmNF7YYr2YzgD6qtM1YdEWNb8UCLMvULPcNGBgDHs
/c5ba4wvZfGAfwLs0XOfPOFY7fdditfn7aVjnIjAHmjsAy5NuHy9FuXySOVGB/9K4X222PUnlHuk
d6tox6Z8t8iwSbmMa9TEe8uwDF+0uJBVhqplsiJ8omOst+7/h3X3KH6odbqtpXPrgIcseGySeEgO
onmWiPxDoYaOWWYM+C6xxk8Z0s2vdgOXtFFjLA5kLgbkjSt8brctDp/zFwMdq9fhlvYMmam3PiSi
EaxMeZJUuYoR3m1bZOBJWsZqYDN2AXX+KSffM22NKp9IiZZH6DP4nCJk+E99aASLciCcv+F2O/2N
TeFqD5Lj17gmKGGA4E0RhkNDjWZaJz2Xtd+Ur9aybBkkHuQNVzR3CeEzxf4+ZQKz3fkUt88FYtDb
3SOnZmVHVr7PZw5Ddd0IGRyLClSYgzE+bGoxuTvTUNrdZb4m/cTFhphi8EFMiEsJZ6v/nh6xMCPH
Oi63lFTgxUxmW7LGrsDDlrCMWjJkj3t/mlna+zwPmKDl8GoTex9vP2nLfitSqgZBNs9G0onjSXcs
d51wz1dJwmWNdKNRJQw2If+q+n3/aFMDpZpNtcpjPTDrYww3YZNqnnIPL/W4xdW4E9rdRWFq17An
ui6XHKOABAia2YKI8UXAi9iFi8R2oXmNhKgOkyUXVMc23X+DCpLeGj6+jouMyE2q+xJrf0/5NkXM
0yhi6pvnyO4LqudePA1DKAY86ezweV4d3naQznFE0aM1GHA4W+wC8X0rijompcrnJlggEcCq4Hwu
asx5gVkE6daOytLbsqKvosIDUk5wJ4cGGtDH+a3A9Gc07JZ5BCvza3COBcULotNkRUpJXduIpdlc
50NtVN1EOGGdVO5KkF7ugInuOmqci6NzXAqQlVWneW6Cd98i0gnilDFNmuxCd/CaCIjpofCtZAYH
7xQvItt53mY+9AuO/MQ6mG1xUhSItYCOzsdDZO7aa+oQzy4CxTPbosAZMRPdeKd8P1kPSIkYelU8
6W7y80wZZMdjJBLMzRkB5XdcbEkjeebEdAjukp5IiEzgmd6PFmDg50czmx7HAbkERaCLycdAkd4i
R0ze9g7XYJr29HNoOgeYyNY8LDJn1KFxPVfZ0dTQbWJnA0OM42Yc8yvlHNPH+XFBgQlj9wuKX17q
7zf4gdCxwklwNupNLvJJr/LVFtKq6nVsaXRZdX+2XoAlEwh5WnKcHFlr2kU79FMIi9TgMIw7jXDT
EHJfrmydR7OYrqj+cj+PoXpH688XYpXv4mqzqm1rciHSK6nJIhiIFjWj1QO1o+umhYAS7IRvJye0
Z6Xk0tNM4Jg70VI+jy9LKbhXprB+tdcMlLxgKm3j0njD+ZqmLPx2yl+U9i8gbiVznbPC8pI+mQAW
xUpNo0F/cSiXv/dQsnw4wcStdoUoeUtrqzkfzbzsX1Ba8pmVmoZF0oj1Baf9EDZ/imceXTy7g9gL
0z+GZ/6YPC610n/yddT0n3+3vP+uNv5zoqQ9zxDvwG6tujXIYw6YfWZY286c7me8RadE9PqTUi0x
TniXj+C9Sa6BeGnoamE/VWE3uAcHtHGcZCqf6oa1fKKbXPXuU3X4Q7lyOUnam9q8hhjsyiYRLFOH
GZn9j/5eOtNqSZiMtdaCDagoaw9sWyRtHAUjp+9Ss/eHR7v0lF8NLkBsJCVwVwkM9Rh0OQ1T/3Xy
zA0ou8ZuzWHEA5HdQmXejx8RlYg3bAB8ieY9nK0M2kkdi6uurdt82J871TvBMRt+EGEi+vmW60uU
vvp84LFVA+xzinp9fsW8db17BMzN2N5CUn3pX603HnyeBNe62XoVQdvNvZKHCNrOsdySDeT6zrAT
WEPdcmCQkzG1nk+YFezPeoxqM59QhEN6xy2/9HGrbbY6HeE1QMDiVIbaSMwXU9KDF7v5Qt0n+V9x
yADaOwXbd9VX6MF7sfm6nNXVWm1B/UaQt8STwcLWeN1evEj8FmcFC9tcGUV/4k5oq9GsYiGs3Fp4
OB+n5G0DU58WYcpj2aHXRsdWSoBIrMKOku4ffYdi8+wiMCzfkRQIicWp/m4GYaLPLUZ6iJcVdRfa
LCCVYmqnFGCZTq5lhc14VHnbhWAUiaoPhwWgIb2OIwNyosrxO8lMQcnwiio3viFmyOZzaEubqU15
k+H1q+7bX7XoId7bVl72xt4O3hJq+GYf9/TwbAfOXyRVAP7AEnjxB8jrYw+6X8A4Ov4krj4hV90V
saks9W5LEEe/hAduSuT4BueLOTIbmQzSnDW5nUrax3BNaYlxpda28GUSAjoG5fS1DpbpYKHxzwTJ
TgSiFuV1Mx17ERFhKTsDxdWAhwYAT//x89W8Y3RxBVo303GY4G3tu+7XImYxOik=
`protect end_protected
