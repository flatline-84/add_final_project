-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PAtHdMJEZw6MJPnIvpnbkXe4EQf5FrQC6qJXSk/xZScSgYwOzBRv9ZGGBi7BoT1aOEEugULWGE6E
cEiTlM1OZWLBQxusFT/vwO3Vt+fWW3x8ow9lSXJtl1Rjd9FyABfR/X8B0QQg+N4PuKoVdMtxjYGc
J1uYsGD5TUq75xI7YghB0LKi7z1+slgzaVsPRWc61/ewzbz1TTIKAX4gGJFPVOm87p8FQ/+ao4Zw
SVdM4HNgCbC7wh73yNSyMXTQR2GVcHdeMt75o8Ge2iPDKlUs0SpD28tZSOtiZwtrDYJLzBpPs5lM
NBWJnMSOkNeqw9npPSH40DW2VA39Xf/Yj3ysMQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3632)
`protect data_block
Df8cPtk+rHOnLXHVoyb9sPHgcgo2RZCd4pHpZajdOPWjrb4Hy60egaID2GRQuclevxY868V6R6LW
vC0R235AHvXzZWhfHzKV55tLHkNuMRYhQoWOrm9IYJ9x3FN2og6GitxoFmyvis4xxsWKcwlq5bL7
hYN90hiLP5e81J3INBnLbadJH+egeb1UM0mJeliu7o0Zd6l7Qsi4gNQRaB/4c/3wE8WsEwrucJ4W
WK6XQZmHO/K/j0ULqIDZESeU2SLJiQfFTI6YnvLNfPNQSzTz5vTd4MGMm3IzGl6x/rq3JmqUrcEW
lN9W19k3BxVPtzxiQSrwdV1miI1vB2Xy2BkTpBqyTWnFYl1TQwqFcxUVaM5yjfVd6A2pUKWiUnDb
h3ar/pMcIRNuCkWpOM/v0nnSpB8zmtAihA3FRZcLQ31qVGvdwLXxkbWLhfODXCBJ7IHJV1jZAsx1
OPTchAX6Ql0Vbk+0ml/sMu5l9garBwgHB4r25HO3XrRG80GeJUrvUIgLm5CdJPrbE4tuqgc2WYZR
hobewf3HelpvX/oASPmBlwX/5o7cckdFGkL6quVxCvbxEpl/if8dumyBh9fd5bPPYgvrG0q+mOcX
Q/5sPhju1NJ4H0AAXn1RYfiY9pwltifGavFSRo3xlWUCWIG8nTnSRFua4GO2Cza+f0xd1Lxfpj3C
j72a2unkRXgXVUVSUhP17Cs+L8bAsxk8HdVBOFrMxZHq6ak9npLK2bM1g+zNchEZ2touv8TEktOV
+/fcGhAnJOOFYwh9NllX3F2oweEVRMu/GK6rH+UiYjHO1TJhajB3Qd4tKLz7+rDC+DwgsTcXHpzV
Na+BTWAXbtO3jRX2q3R943b5sMryZCaGOzHJh+D+aEUB1YE+zzzbrmbfbxx8jAhkW8OsuqWWIk6U
KjEIK4Zo8HRsraKkT5oAFeWTLv7eWrfZ0NVvqZqjEmOWwZwKastHih6ninULLOT+QkQ4zBBG5l3n
5weoguUx72ewMQR0Lja5isz6HCF/Tt4FJOnu2FA6n3O7vux5e1zv6OIJW7y37/dL6IJi9Ca3i4Yi
Le9nx7+0+jIgOk4AaVMnr1cbSQ7YjUyIFdgRuSzN3ZDR82Eq4A6oDWfFFzaJPA1/oEajGpz+8GNL
ko3DF7bc1RcfhHyWZEiyqS0uR1CzctJKFRNNDYOLkKA+SGORPnMlEPo4JrTDzhlMzj7F4juJ0VEi
Db07lD2ogzMrn1hE7+qTw/uU/CiZKLCtKhCsNHk44JS+yjmF4EN4kRHyO3dJSBVClTER9R8LLPX/
G/Z8MpkhDMJQCGl9Bi/g91N5DvbbCmE/Y2EphElZGvMRbJ1QXhzsU3W6GXQ7vMghm8EP+QwBGNrf
TY+u5kgsmrbI+MRuJGhs5e4n8K4xfq/u0/X+rP8ZhV8l3wfg9PtlKqLPlmXkDLHcx7h5H8isqQFD
g4jMbezxQNt0qxEjtsX8sTCP0Jz52y0IqA3s+Kr/5VN1heKtseLTvXg8uYCP+V3sIvxurl+67fqC
BG6wtGFgOT5T4RhxYw4lt3fzlOAJTHQh9oUvICe5MQA2/iAYm2ZcVIZt/J6AcQk8Y8KlV6UIYI3e
oDPErMG7PSzHd80lMttySaB/BacpgNyp119AVSXPUpRYqA+Jv9ZPaJXikVoIB98R2mN3P5bARn8w
VU58Icd5v/HcmKbFMDrKFq5YEE1BUVDydKTsry2I09xG3IYk9BP4Ifk1opE6G5ohBVWPrvKjIJaC
NFGi3wYXjuxy6LdamLY8rnT5Mem0BGQU2S0dTMAsCSBIB6Pd7w61CMhojFrjCmoZXhddyA2FwTIF
u5OQOpB2HnRZVpMGg725d1PvNV5bWC13Bw9TSKKVgjEmKqg0B4/HCW/ko7FfU1qSS7vvNfu+CXov
3lI1pMTC9/CZoCC0czTl3pUG374EOyupmY3Q7y/veMYuXY5S0uBbcJphnWJTQAIeZ3wVZ/d4TGRF
q+ni5YUnKwHkQBVCaD9DbUPLN2GimBgIddIppjxTX7LvAdeocQK6fzHSIms/Jfywg9RNvoa/E61E
uAgCr8sfJdQEA+MHYOli1QjNxUKIBlO1lqPu/GawehA/5qsjFPybszq91g/nNfeN21UBspCWarZD
TxZE3XPAGb3qNKeF+nbiMJqJB7i8eE/lvw8tKWb4zu67p0BCltfOHNt33K4J0nxmBnqnDco+/qEH
VHIRO/mAaj/v3dT6be/gytMS0Ip1pyGHuy4XBG6EJL50WJy/ghValDh4l+DgplBuTMMkX/F5Hv1d
12HCZTNJIM8ylC2uTaFhHQ/Ubi3yN9OUTGS9QD3rOuZW42Mmvq4wmJfwvzOz0XlonT/lMKIcgndX
pmD7sRPlqpU2YE3aIXRBjtKKBla/A9GVqX6yyCc6AdrA+VhEpwwvFjl5UUYSp0kQ4W56jrk64SPn
LeSEDG5ur6G7FYmuhfinZ1eVQY84t+tVHUnN3UgdTU/Hw3dqLaUiMad9c22SZD9HHvZSmImP8zWJ
eZfoXR59El4hveaB89xGHLb+MewoQsMQnz9I/KCVzJ0nBn5qkMbz1OX6mvBoTQPw0sALr/M7l6Xj
Haj4JOIr1/OW3ckxa1/iJVZMutYiZW3AhwNVYsgn7AB+TUpYSWQGqcoFDTN5KBSqZXkaLQxC/JWM
+lQtiK97FytvPF+7gAI0PngmgH6JYIYNTg9vskQrZD0+BNoDfjbPcJzHQ2TVsIr60oytw/twZhrG
I1zMnTv7H/LQooJfU1rOYa6CWXt9Mkd2wMLwYUk0HnQl+u12khoQ048xec+bA9TCttOVjTljkP/4
6vCYNzko8JUhVhcOHcuSLjybrlsuqlrWxCLIC9QOhre/xoxtUP+ICJjAL45tAMgO4jwpC2OUzNHY
FKniDBV9G3dDG8I6ifiZpvnUwbQn3x7kTzQImK0rzFKRrLZ3nhTUbhSEi4Og5QjRP4I48WPDEZ+o
Hs8dk+kRV5Lq/mLmLq8eiBNG//UMto4DigBZAtWfOXNpddqzGAvJYFVCdIMJAuvTA6bphu7oqgw0
jzMASzJAJbk7Gyna3jJokbwkAd18QD4Qyr64ghkTwgYXhlrMd0iw1TUqCU5Zti8g6996rSjYQI+j
p5AGVY5W6MWnJRCmIdurKq09Tor0Maqm+Ab9DzD13jzIUekQZHLZxmgTq7SryvbTDp2Zc/4dJlVl
8o9J0RhT59N+OPcAAQtgeRAwvdCLKvBN3W+e0FXCur5KEcocIMvIXyM+ubCfw3UzujAkgiX/WqTQ
Rw2NLM1vscA3mWkaIWv1cgIK3w/Ty17HaWt3AxI0eRCToSaAvR6EEnaSmgPlNorkLUoZ8mJPU/Ml
qnsuu8GDTajLoWzDB7vG4i6vzKmyBOKBf0fF+eGhbZmZX64xs3QGCKy2mgQB6a9lTrP1lpJ4bXVu
SI5hfMEUOXQJ0cYkLX4e3+uaaZyCio6yfHN5Xy2CrtzRwsC0YKnEwzvtO2A2fHGb2L6vghDw0bBw
ZzV0VOms2t7PVjHGmB+CHrhk8MuZ2Tfl72N/6ACqY/BTsydFVtbqIR4PzckatCl/Ap7ffh0z8ai4
grbKPlwZeiaHzCe54fU5m5eXfvN58eR5cY+XO7xZGDgqs5wDbLayX+I6dTtbKur48FYLMJSxmn69
u2jzmY9gYi30lehzksrpmrXmaWByAVBrszRxeMANI+hdCw39uredUIMHuPg5fUiH+S6hkHtZZI6E
guUi/WQr2EoSkrn6Q/kYGoKt4PyianOqeKfGb1e4iNl+OFft7CjHm/ohqy6rAisvvDhhj/j7c022
kW4XtucgrkhylfIdN/KpLs/fd75LrZuuKEVordXjoMno918wPrBIQPPoTW8Bjy9Hk4Db4VsbLUX5
97rPDqn95WM1ODBfcE4ROuUx+npd4W+1ZXRvhA3ioXwGqD2WHxenMHp3auiw9BylZo7ZCS6+MaEA
wtIc9uiPK61sGYfkWKXk9VCRxnf0QXAXF/aFj9zyMK1XpE1kWnijSzW9+SgihhdTYsyXwnL6fMfv
PiYXOJ21BnFV91cfm/WCN9tBOPceS8VQFDafp9wYD2En6aCU1eGMR1DSUZlZyV3s3wFv8l9DpWay
H/Lm3FNkv2+kD2gBRy7CgOyuJbcvg0tlDhEyk+dJv65xqtt/6XIvOY6rpBZg6bQtcibpr9iYv4wB
3V1/cf6eTsfKhK9ePrPyCGooscKyzFfR5nGnbfGZvZTiEAIjg+hNNfCpzOWuX076SmVWkI2CSLz/
lDzv/koEyzLYbgQ/qYcV+2Jffw8bgaezyZNSfIdA2PuiqDtJrxoZna4I9P8JQtfpAy3fuGtHq1iQ
4uvep3qnzQbd+NRsMmoiJKp271cfQh6nk5oy20H7NOr3W3PsuAdHuiF2JryJPUkxCoENuI674KxI
tbU/UY8FCFTKiUBOaesFZKft4BtPgkvakOmWNYtH6WxKyb5iuohFtljC8LuGCBu1ckVSsRB+ipzS
eZVDCfzFxgW4k7eMgtmnO9pAN2AWIIK7UKVxsjVXlOy5lryS/5S7MWwxLDDTSxwF48o5b3rxS9Ww
XWexzubJWJdEfPoPIoa8MGGHZw4SxmkDpyrB9zoupRDrbgrC7YD5e6m208fUNoOjmKpXLigv1kGs
zrzvwCQcy1t7qz3u8yiGt2336pfMmP+U30p7UNxXLEV+JOzF+2Qpo1I/0gueTkOofES7rIIu7ECN
1WYfaim4mUYYGNEcp1Qnon2Lj1Gj6XnJIYBxF828TVn/zC7Kjpqhf5u+e9wUJSdAEGoFpSm4NX7r
G6lxhGf5M0znbH2YEEZl9aXrd533i/zw09L9oEU7PWbCP2S8NcXRsVc=
`protect end_protected
