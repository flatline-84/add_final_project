-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
d+bX5b0Mt25AnIw1nGQOW6+BfU+mfUgiRNMgmWY5uN7joCrqy1Y16JiU4hqL9begfqx9cnR/MJN5
tA6DSmzqxixsLzybpzffvgJzsZj2N0ygK6kjdIHEKtif0Z2C3kigxdmVtR5v606nUwhCV31RsY4X
FLCyRjlvzUM9b1zP9RULXwjexv1SXkaRWspMZeyQzDHVeggQtGDCM6DoUvLIWrOR1aAg46ADiiuq
U5wWzM7jYIIuGPxIgCRUGg/k3v7abcXfWBr9X/PWk7TPLJEaQuoPTKhXczh5JuGwHi+I8vQKlTEI
zJ6f28dz5OvX5vlEIpVLMqidjrq/FYDGT1kfRw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28736)
`protect data_block
0KgHD5UrReihcqxXK2C4j3bxTSrnPhsA/cXy1mCXDWSLYxiqxSp5x4cLrxt6zaKfV68kChN+uwGl
S+zPM8D4fcwP0xXDRth1S/9KhgIPOMGE2F4KUzVpBvHdZO5eVqxl/QYjDMDL4TshZWOU4SiUsuQm
J6Ie2pMcRSlp+1CCrfuSBbfTirBYHwQmS3MCmqaLtyLisUO+rpMnd2wT6VBUonK8RIYxhTWY2KtO
RNXA1Rm3smBTqyqqO0wI6cs9i3Q9CA7gkFdgcL5TnIOPYotUw5oG2Z8VSUhBKt51lroWGzySRkK+
LJGSfT93zgfi11EGUeY2jbtqQeoFun1hu7o6ZahCSXTGuoT/q7lOX3fbdDoEBOpa/FGZV85YNSkx
QGKr2sfM17L7U2fgSWn5RTiR24rVWLNHBVmi3cDolBSvd7oF7b4er+Uhp7SOZ8dTG+Jx1jaiIaeE
/NuZjh+uuJjIRnmGGAUDr42dYlNhYlX12RshXj7iJ055hl46IwA7MjfqVLXthrQ0B6ZyVqiSrCmQ
kHhSDIWjpcZgJqMTsLKX2uLcDXmrG9mA+MhH8JpRqKc2mpkUAREOQJu1t3LplrM0jGQvbiURvDwD
EmCRCsDEU5SZrUrcZSOXeiFtakbGJgB75Ec81ka/KD3cHCV/9ZqwamVAKF2bgPEcMeEzzf4jXyZY
1Ne0tgtCcAbYQjndNHLCNNPm1i5kAuKNdeMZfR5B4mbK48AWzgwnGTqyGezg1+HHkf2SBaZNQXMP
QV8x7Awp8IcPb6zw3p8gwvdlmJI9FjZpybJXJgARSKiH1JEFz56YsyYv9yBJRQY0Lgspu9C/qUpZ
LyFiAEaNd93vdtZFdu/QNzLb827eO/U/uBw3nMH3KkjPafmmJLARYxDALCD6V7E/D/r5GlBAkeCI
V9m2VQWd210ly+LCtoR6VlerwN97OApjfoui02fmtco8RrXPFimCf9tmun1D+ExQGuy4++x6NLKX
IeOBZlu6w4jJcZtN9JoefaMG/Tt6K3UME6dpKqO3OygnxrEum8azfVF5TXU2SaXpmgnrsgiRd+u3
C+ag4T/l/VMjqRv2ntMCtiNsCxAHR650kA07wL3tpjEnCGEumnOxL5ZcH9Ifo4iyiR5XV6z9vtQn
LGnk19lYb1T2xztrTnTow6vrminaW4RP16SJoPygCF1W7IeoFm2A3Sp9eKHGqMTTQAETxXs/3Tl7
Do0DUhdw8Wf/9hrvIDEpK1Y0jpsxS2flLlosg/1YE7Qi/QKolsH1ZvU2lAUAboMDWoTHfeEfyxz1
b4mDh1EjkyOqNZBEpMXLJo0IgTSx8QPJfF8GvPw5FpYPWtlUCLtWnQyNObYQa5ws89cfsN7g2ANl
tvjn+rdYDaukaN113muRL+PPPAGcOTrxQTa+mZigNFMGwDjRTvYedZAunDr0RhCUR8Kx/OrN9oZp
ETLM9QfcajGMDb7ZbL7qURXfAhq1AoPPoDqWeVZD8mThRx8MfyfF881Z2AfQTASmFN/Y5Y6xC3HJ
3qsXKfkewgnMVdi5/8vZvcDsdP3Mgb4RTAD0bxeZtuZlhNvWvNlnZAOVCW6u2MGSrRiVSOMjEaA1
u9KgrOoyI4y81zRMvXsmXbc7K+w/9QZJtBP0C5kbBGm3T5lpVfbQSg37OnxaYoFfLpCj3ErZHMWZ
CvarVigeH5JO4uBhV7EwRkrNGZshVLlIeFyLBuNtqk8AX+3sNeqCQatl8WeIn/QUdSpPmR0rEea7
ea2aSegmByC2MM2VWg2h0kNbKD0XjneD1KcexdR0DPcGjJo/pPdM9tuKey0JIrIcVj6SXZanszgu
gWaTpd97absoHRG+xSJVpjuzPUogWAsBKdjal7VVyjpxMz/6ay/uEdRTDbJKS+CD29ON7pm1Tw/L
vslsQZiBw3RPe2NSXHqqWHHxuEDpaFfEWGcyq/dEY1J2m+Lu8yiFwJQr4pR95sROLBCDh66a29bO
uRJTvVRV62ETEb4ouSdna+q/d1QETGv5iJlsbZ0GCWvtJtf7LLFFZFfiY/zgz+nkZ/wn8C1OOn0M
wD3qCYl6wn7Qr3BcfSdRi2U0aR72YG8PFB5crVcGKeH2wtrmj+9EucFfMSexmJGcDB8FNpIQBeZx
VIrl0bgqoXv/A9uiOnFYKQiZoGLhwI/Avqa3wVwqd08Si66CiwrB+Em05QV9wo1WuWPcfqAQTQp3
BjvBnnvswLz+SaqmJZHJGR5ZAQoTC7XQwQ51qOHxjW7IwQtE9Mq63qlROOVNs4fwdpAXaSE/Oj2Q
q553pMuXphNKSHDI2BH1br1aoPfcBBcs7CIwLwu0//DpErp9HYMsMI4qJP9VFki0TC0HK1LToRNg
mzube7CLEo5ptZfO2O+VeE1Wm6TeXpM1Pdlo4Mj29g1/uhymb5r03Ut9LH19B14ZxtueOIOcCNXW
HRYOa149UWSiiO7lR8F4qtGwEm1asBNPHzGzMuV2Om1w/iqkB1Cnm6Yqj1cdsohSrcq0RH1ei4Wz
VFb1doZC4+hWMeNV9X2HDqtP1dG0TU8tffPfHqlAps4ZZ0hPu6w77ArORty/BNESGVxvPKG4q5/P
4qiQOaVXmc/ZZjoD40SKtkGCra+7dL12XWLHhshskh/SHn//QKqT0kxBJIMwHULAFjrhL7dLSXdE
iqkkznvEkGDqWyx8DzukZYnpiaT7KRQ4jTKAUuSVojI9C552X67DSEnpq/6Icc73n/aD6mAabk2c
rblz6ODRRPKCcCI6jBOkXarwTXfvYk+QIatVp25o0m+X5PE7ALY5E1uYVdtbxFHdrtWKY+7nKtkw
CSEvLJJ7MVjMfF1XAE+n4X3o5GbOG5y5AaRgXmNrb2ksyi3ClcDLqHkOwQzvXgwOCaUpFrF7DzeX
MpymffuogO3do09YSsAoQ6mmircd05sMdHfqNk+b8oh87W5JOPk3he7rDaW/l4WuKJcyQEe3NmWx
1MvnZRCs5yU/eQB7xQcDxIlEF45QjgAXIKatIFVdQgd4f4Fv1RBankVy24hlqwtum14W/dt1rwZp
LzUz8LgOz+OC8veOzx1pNwWKZ5wjdtH5i7hvxWVEnOuCCwGO2hkOlishshmWvLEggWFnkFKoPNUp
HNY61PljZpWWDS8d3jMclLVq28MY4Qdt/T6VViY8xrNP5mInCVDrm65NqnfT2yGL8D57u6LbXgNA
VW3tRBDjUFqUYe06vsWEgbJjO6Npk8gZN4jCmdHJl1U5UDGAchjAc017qZutHAjcKXMXW2R+dvjh
a9D05AfOmpjnhjGu2ABWDlRStY9TWSrTlHkXJ3aehPMeY6kZSKsRkJQQVKI4Ck2fNwomheOb8IC+
4Q2JQ+VnaWNJF8V2EkxydDdXThVq+/G1BxoVcVuYdH4dwc2COC3zGGA6fb09j7njzb0Xor05opz4
lZOI+mgGBJ8bL0XyqEz2OnsA+9m1B2hm0a0/CEqqxQLU2d1jGgBqFUyUyib8VdEk6OpjtfPlVafE
L1Bmvrx7/Q7Iha8SVbv+rv0fyj7Wl15s18LDboE1alapAQCumGkr6HoYEdks7hU4MQdoX1c2V29l
XYKjyNL8Z2iFspYCc72RraF1us0ydN15QzLM0txF5q0JTrBxFdqiVh45028dlLtCWU8F7oNzEDMl
7RbnWUkWpZPuHtWw6kIOUmNpEGsRQo7/8IOkMbaB81QwEKh6MixbLRg1UScB7S+NI5suG3DyxOuE
6O6VOPKPfg70pMxH+XOq14aLZcVqNRNPgpPkTOEdiRKrI5MEHIjtbIDz6b5RKj3+2mlJILfSoS4+
/jOuXhrww2Lh51ud8Jd3nyquHX65OYiS4hkwO+p+zM8iRMbpFvFkzvv74Os/J6Zw0uM3fbCaTV+V
nFRe5c6HLRkBN/HLS5WZoXqfZqRP1UCCJiJRynGn0RfA36OQ0fX5nWwtQNZnVyEoReh39h6pyWgm
xh5GtDC/pe14SDzFTw0yBnZAZ2WUXr4zNJhQJ72p0WmzftcjDU3dQGOtw9KuAgLcq0MxNt/L1pRa
1fQaE2uc/TtuqpRJH8cf40LMzl1f9/PAVtqTLVvyrfhlHcYPNWgudbIV19FD5zND86mHk9gmGTQ6
QariAAC+8ToXuK9SEavb2hGFS3a7XuljpUPlEeAV03JOj1B89DKMniCkbWWkGkg+Dtk6hYlAER6V
zW7GDC0mxZ3Hq6t0a6aPzwTyd+7PAyNvzKsIU7jJK/cMWYDsc2R9gYt10a3wmy3dO3f5lh8n5qYN
klIoWopmPHW8RjDaiDXLGkS2P9eHK0C1hBf7KwP2uGyPVacxfflMlD2fdVoUYp0NX/BQgpkpjdx0
DWkbpuZqRs/0jlKfcYfPbWgb1RdSbL2XXIAkWRBGqco39d2fsfe2TxZC/vEVE6Yd0gV99Dwy/E7O
rdQWRaILVnBBQg+vY61wt7BHD2XWNMmfuQDRZhgISJICCqyTlgwFEyj1B4iS2+sMesjcxUee5vpA
y1Ql/4gdWlAf/PStajnVywb93+EXHPzZ4e9wjvaIRE13/d48JAlQrJ5oqatyTYY5vsJ5dObY6uhN
/RHjqG4bXvwJvthu/UsaW66a58EmahbW3neP3r3HyPRimwbbpoDDb6oF5L27J/G9zUIn2AfHz2dm
zJAwQPcpfut2YniEpbqpRsERLto4kkbrvyza8O7a/5849g6I1tV3+wHOu6mo9qGwHk3ky6dKzSsY
UAMfeF2bF7UTUtVOkxfKz3zQN9Q5LTo7lHMnZ3BJKb+Wmep6fab5ZxsRTPEP3tJOTtpEbbpHcU+/
zIIcxzJWoIze2mb1zIRzg9+/dkrgSBGtMdERKSFJiP1jInVgupWrkd+zIlI1Zr/KDRc46+UIV0fM
LU4IVyHkbF0QdRK6tviLRGkkInPJaTWTxBLSabcjyPVh6L0Q82gnEOIn58LcYZMzx7oZB2qHLWp5
b8x6d0lzbXWpuc41mwKKNmYH/KKV5CVhiZO4hjeWToMfOkCLRVFQmUknlGwu3vpjO8kAlJ6OsjwQ
G2cnA9N4JRpZE8L6jd854wQeOI4NPCRkxZQaCViVcn1OVmpIyQIdYDEJpRM8j4ur5D6ai0/fb/R0
YATSdQuQewYtbw+Tjc4XU96bhCW7EcZguCP3KP591/rWI951dcIuxNIuZvHuUvLdJIAOw4HDDyxk
9HuraGWpzXfMTFMh/QXQ0Wo2mZSbINm8YAOFC68rAmiv32XGlmrs3ci70z+JD8mr+vVND3bYjKbV
Q1uPEeq4Jth8p9CPP5foYP6UcUJsbYFS/P8+ZzuJwhqweXtyuzkdiLCN0DVzF0zBX4zOHPBvk9Z2
+p7w20x19nrqhtA/ibEHoWkur6fn6BN6G8YL5dYQuvyDFcEP37rV3hyuRam3n2bH7tIhBJVXfSCc
ozzhqP6Xr6aNLx0WeiEtdTpFpOQQoBLFPUXSkMiVzodc2/5dbuew9qwDGiJ2vZ4fZbdFFYnG7Eyf
79P9U5FtkKoufn8XARwdAJqGj4tCoKSBQKqyrOZTrM/eQhvHtUCJdfVcR3JqcR8yAALwfsySW+4p
zKNmvN22aySbOlZwrNVzFPJR52QFYVs9LnYT7S5Dmh/d7ZcWoFWn1ldnbOacy1bj4p17mJg1NUDW
pvbvvSiBpjia4yeCYil481L7X+YmK+8qXPqNo0iGX51RutH98VjmnmKHHl99DP8y595O7c6kuWpY
XYPgjwvmo+3IRT5cCoOCWk7iLnA+jmj07gNj7fRZWUygVcTdatcNmBChiNRVd7JQgWujKspS5VJu
fErbcWyqE4ooIQSG4dgE0LJl7XjrHvxgD7k/8cs0An6L2A+cX07UyPn8TWV+QwOWjvcp4LpQdT1n
WWpsyHn76TBgZs1fZm5fNJGuDOKAhkrKag/0MzRqStn2mCCd7I6cybeZ4vNCaareWrelfqS5DwHD
K9iFvHX21WRJQjaLU2b8x0CbfMiwGfEbQ0hOuVFx9hS80OnQA1erLN5WlXvsN86bnol70/t9Okl5
cOXjQ24dGoGSkpraCLk7ysBPxSUp8zXRuVGXTNPLaWkJOQXpcYe5xfnUs+duA/ex14967rdYiBZW
8T77kRPfb/cDBZQ6Lel1tM+SzRiZKb+76C8RWx/IikXmJIzCJKgbrn4GmYYp98p8v6Ba4Ps40cZK
HkaSx7mXEi4pbbyKLQCmsfdZD1BRE1v0WAg/VBk2V03s94nFExwpb3Vl7Zbnhid2+S8qfLpJpP/F
aQN0VkU0XSdPGzV5cKdigVzIrJ1Ew1NgNdqKyBkcjd2f8XD4HH9y6BxLgGZDGBI1pFY+EgbnEeWT
J+syYlCy9N0baCbq5yEQCZYyy7AcI/O+8toLuksBQVb/gkqZY4AC1mwkEjKr004q8A0AxogM/z3P
rZ+5jk3w/BC60nMyNFFzJ2OMls+lbjHUONy7J86cZ+IXU2Rx/vxvGyxqxGW0CR4GiAAP+5I10YFu
UJw+aBZsXjzXR3d7d2NNHJy8qmVi/oOg2Vq5zMLA3nZNdIkOqduFLzb2js5OHR0XMJxUUMjbqGYg
eFCIDtlLN5f0Kq+Wqq/l2NXjbkFb3Ofpc14QrSWUOd5Yc5+5r6M70/fy1VWTt6BrRatalQilCnMl
7yjCVN3oj0mHZF4exey0rYZh568u7oyAuiCsmKzr2bRc2XZ1IumVV/yBm8EkG6DQj/5b+UjBab17
pk6tvxjH2n6Cjdi73ifCLsl0e+Yu7a6LJB9JN3cH/sBzgFzC3ivRATXVqIlYLFXSZ3JARxw2KgCB
EL6yam/GqMVrDP+yOmOixcj/JPy/NrTNoG3VTZqtD1zp9raLmfCd5SazskcSe9fdwyzQZGGjULWE
PKaoQa8cS/CIcK80pMgyombqfOSx2a4F1DsO3FWmUNKOe4u/vK833lLdwnhz9t7iNlTDc5z/mfZE
1DhBC0vyIhcDqGINX7/UGR2ITnHUG7+u2m/x/Oeib/kiBgY80YnQo1+jeO23fhzQ+fhA+fqbzRue
b3/ursi8OwQHE6292xrzz7tMb2Pus9VO4QbliZLFyItL5MT3QIWHuspYE7ZRxODb4+IS7IyrFWiO
q0mfFiDz0j31ab6y1tcup7o1fLKnyD+Ecy7fICW5MbN3lvcgTv8pGugV5Q5ujtTDp5AS9W2UpyYU
Hzi9767CD9Pq4Dr4Uss1hettnwIETH7LgEI07LXQ6dgAqpGtSxOoJrVYWHwGTApVRpt69mr7Li5m
eyZ/h1WgmgllnpT7ws+UmHcx0+QSa4FcKjosgXwA4Cfdx9AEAht0sM+hi4KntO16gNzwP+rQhOKF
vgbdvOVOCsSyLqny8T/GS0P2X20DwUmTXF+tmCTzMqVLdcEk8o+u8VpF/AsT/3gSzkmuJwaloKux
JmoAwe29FYxx7ET2cFEBywaGe9JcvS5AxWjN+hqOC3XHLLV/E/oHqud4RmmWYORPU2Qg9Z1aoU24
pGDazTihRy1z6UsCNZnoixpZ435jN1pr6b+Dg7qyHAx3BIzidsQ2HILi99cGGHx2PN99f2cHSJBk
GqjOnugGOvFUABT5xfzVoJ9R8p44Os4w7OBp+fqw+SZBxaoeuVydEqVeBRWzq/UgiDajAu159KHD
IghdYpavxqCcRSD5GrPHe/vZRlL7ivLOvgJ/19EU3jN5igK9uH+tPO2O1fQYQQEHadMjXmGbvnfo
tIIBop5cyCy2Hgpx0VnlfE/uL7VEkbIaKdfg23JlWHWkOtmsSJaSNJIfHJyVGaD6trsW1OddjEKO
+v+HHFgbiPrObTprq4F8w91ngWiLc5fUsRbphcBlqtc3JkjAHTxfzr7Zsw8MYILwU4Fvpz5xXiXu
f2rjwjtl2hm35lO34MQWhLZoL+aOjo0afeltISul92KULPWUYgQ0uve/dnxfdIYbOH+0w5IMc2YI
7USblO61jfA5ZHBvHal1jzZkrX1N6RfAGkKAu75FvMqTN6Br7wrt67dQuOmQGafCmNxAhR1+hwQu
5dOuBrasZ8KXD8rpTaZ2q6pnW/QwYjUt/LCg4jXkwAuIiXhEj9DqGKUhLX0uLnXy9yiWZfvm9uyD
i7EcvZpTvhiuy3hT22D1FoV3pn1qx5vfEazepB4Pdpqzl8lRRwFQ0gSzpIlQEcQfPeuG/bMBpOKN
A7ZawqM5tU3rfx7wpNBXB1jXYcPYSoIbkvC+XLV34CvFnWd2qmJMRYMG1PphlxS3NLkONbpM7FsZ
F5UUKpk/O+K7c+LZFRu4ZNgvMFAZjMGQfnBoe3wSK272urju8WZiimyV+irqNr5KPAeKJlCj5/0b
njcB7rynX40es7SQhWbPoDuPI4lRwMa4UfZQcl766jAVzUWWQE/UyfxK0KVNgbxiXxh8qAqqIpib
sBpHBhwRpmtXvVrcvpG58fpm0yGzW77b916E5F1XTKpeZGmC2Lece5godJm2wCUsHADrZYtbirMy
SbUjaU6QHbvkcn90jYunNKRS16Z+DOoBzG2ajVIBl8b70JZ6npu6kJCOd3ZI7sM8i0QeohEK56Wy
Axts1O7YmrrcHPn8hGslTsUkjcV6ag4tFTQnNfSCJ95hLN4HcwbdrL/iYNlbIDwVTM8W+b4hnEEL
2G6wxZ7np+nI8f2dcqwMVTRJVRZ8KEPt6+f/fME7D8rI+iUFKI4nTLpn5bgvo3AThpt9dX2xjlk2
rSyeoI7xYSOYzglo4OlsAxh7f/rDmpO+RMxMHA975EaahqOhND/T43uNvOU2d7aVUPSKPl8Iki6+
TMFsG5i0AXGM5nQqu53aHXjegsd+gL5ybmbiAgisXVgQaHMbBX3U0Hp4NthxyBJEUeAduB0v/J3N
z1H72WbTUz8Nigm7gkWfmaWp1vKFb9JHM8pLKpcXBLh+gdcXlyIj/HCnTkyCmklaTMcMxIUokEfE
usWqpeo8UwMelrt+sl5zUFUdIFxJIDvnP7ka6BsMhinTGw7yrq0CyCL/JPjE2lOAzskQi4qKZuxk
jkCqAHgGuNWFT8p2KG8eER0Jv1JZ1Ojq4WnjglPPvMLMuM9OFnxe7iHN4kaLHX3pdfUm1ip5Mr1I
gUW2+xogIf9AYfgtJR6jrBW8zdvtKC57NZT+1znVkMr996prHzecQPfRJS4aaFfE+in8KEz6v8sC
HDkTy+Rd8RWo01kj/iursl/TH3IWHOg/Ri+Zm2JZq4sM8heWaTSwBLQ1Cmh2Dtacm7/34iWoxKCv
LCvM2wPco0ltqc3HWO8CaPAfXEGSsqms/MI5HANzxjiZva0YyT3uuCdUzz8cGw6N6tyl16pkdMRP
c5C1+i8KBIoZjmnDMh/+CUxvkJoZHCwGt5GlAWzdS3Ymnv88Iv8tOHL368w54L8PbS6vrYpy7N4h
SbKtc0MmS8qSBT9xzLPVw74T0SO5rCFZhUrCZgnXxrhT5c7SLWV0I2zWHDZnxq0AjUOrK4ZpGdBZ
LOrQT5498sezaJ7yoAGhuLqpcI0FtCw43qjOnuOxNnn8il05VEOXCtTdBCBP4FKoIeBIi7diMGY+
gsC8sRhE8R4ad5YUorVgzejkHizTC8AOoIYJQO1RxsjMFpCd3VSYbcitFjpB/5fi6B5xsPl/sL2+
HTTndoaHcLZPfNfpa/xFHEY9nXyQMUSBnId5aqE501zxMaO/fuCyqbvwfqLcM6qrsqMx26N3DC3+
JnfrU9jAhxQtRkOj3qVxmXLGl7uSC1mIa7bJO1jFSU5NsO4WwUbVs3OnchP49OFsdxQGo5mw0T9L
7aXfWZ8KTEI3OmfXDQtdnSAY1aPBmEQXVQTW7Iweg7VBhmv07tDbY8J4pTn0+Pj3T2eIaoO3OPOm
UlKJy8vRIptr2oJJP/CaPjnIFljYUa4ypa7rVezlHbmwvCAFU5ZUSXez3i5kv29l3S7UFD6zwMja
HirArLJlXS3DizsCOaEpXYj2ixYFwPb7KABE2WmcgaFkOsuAJnxLtvw3+uj/1C1bDr+FOO+TYDIs
/OmeOVdI0xTQRy/Ax1JQJWCIq23uk4lArl2JXnkUANWudSYOfjNX2TxfcIZdtuHpaBmnpfEIX/J2
qM3xFy4bLkloADDFY7IHc/qFWPaIZ+LbdWsQ6Yy0FlkTn4EQyPoI9QVqnP+8g0qVX27PS6MPS306
TLvLH4WwjhsceRSN4+mdDp1D5CzOgTH3wx5Z5L8bVj3sGRdXiMh6WCYS3W65h+GkoYhMBcjVfFVp
ezaIz9ZvAok0ocLHNtQNMaz1ZoPGO5zbG9Yxa0mbbVdns8RyE6HA9j7eZQ0PMEj5OHlrJhIqoaIX
v262qnCnoS7OMBbtU499/TdfS5TqS7avzG2WGkv1TLS0surNxLNFkg8Thih+tOfL4aopbWw+ZA/1
k0kIv6pfhZdWWFqOmM6ZU1yImzdrZm1IpLNaFP3ihnHmMBd4sOsZVs/4ZWjbM+h6kLNRJiuK06KS
iM/R1zOEGn6nBr/3T2FWVbgTx0W/xjGeczMqM/G1K0wE8utTzy8iksD5PNF9rNLEMcmvodQSQAJR
DPZezypWQiK7DZQmxIQaeAEz2vFm5pJ9Cxdduk0JTPkwYZQ4J4+7kVsAUr0l5QjSAwISqP2KECMV
BxZ0dRLkP8yBh7dA7zp7DZvXiuscRByQgS2BlFI2b/WKLVhMxJv75PdxmrfK07/YUdZoDYz9U3lO
/spYA4NxCuzoRD7Tjadt7u9L4h/RW4S/Nd9NThOBXX9/Yk6QtW9frtstyFHTY/ptLYAlFp8ZeImB
LvWJQ9HbSdui61o1JxNOFjPlTyaEvN9VfZbEaCD7/1FuIr50Ky4x23/jXmXsNk7fSXdXIKw+iueN
AZcCA6vDFP0HxtVT1YubqbaBXB2OMaZAmc9IUDOJAIt9smWM3fby6zigkUNDMXvaSX6Y0yWiM4fP
csUPqV+ilAaVWa9xOL0bdKCVmfGjmcBo/RS75kya8tKRjWXmxdtzQDtDBXtUP7qylr/b5cUf4RIc
qqk/NJZptMLPM+vxxGWUniphO85Raoj7jD38P3vvQPA+OAW13NCWNYMEGMraVCVcymIIFaW4h8WZ
Vzj35GIGee3KOVZ9oFteUMdGAfnceCTndVHCKitQ283txHz2COSyuSpdCGmffeBFcZSfd2rb1zfW
gn9igI2eH7TTUQDcsY7CRYRtiOA8xP3dqBj0itVG5LgnkbLzXNI5EheYJQyjOU7WlPyInFBPAtH/
KU6SpC4fAwXDKUAV6CKcE+VJ6pFDxqbBwtjxYv8mC1lb9bRJXfNJdwixvZpsKXo/E5Tlo1Ljb/xn
df6iGxunfD4eT04UpNUKQexLsduPwIyr0tPyWwEGIk2lSdzkgzoqU0zKYbIEQVpUyATMVEgAuZml
MNZ6Bp3SYVRZAjQFkQ0m8hveNKFy8Hz9vDfsy1K688cjwVTGsm9Qj4cU+jpMOG68FTtmRXbUwZt/
k+wK6DwqvfeQX4zMmhsMWCz5jOlMZEsmzaArg0CPoRm8J60MuJRBjH+8cY0yGoosx+X7bPgL4Vcw
14CPxNCFE/GRmqv36sjW+2lh+K/k8OBLAI/MnmVGnxCaRO//YWac3cZsQvOFJsaudo17R76qRYyG
/IazyUJDWI7/N3Et7wszBmtiEnMD2bEZU8yDdq/aOwDr88UDFT5CnP2TeEVSK+lx4lQbCynoQZJr
UFriJv4f/g96cLQjvNyw4nrtGeWusgUtHd5DVhc5WZESQiYGn2HdkfiDXcb6dOwb8dbiLL7oJ9Ad
3Dm4H7PyqJfnZB/l13flZ/snUQ3Bnf80rg+4eMaTqUG+dpTaJFoyWsVc1s1BvvMb6cQLT+FJklZZ
/FCBDHyjTVJ+QFUPVfztEwOFvTz6n4SLtAkaKjf6sGjO7hDxSsR6CXWPmDWwhCseRFFVqf/MFzPz
U0lh/e2fd928e/6j7lutzOZD93WcUyT0PniFH2xlHo/HR4OGR6Glf/PB5chqWjIt2X/+DZWpE7dE
/KoiZMnDpb5PzjvhoY3jjit5/JtfKXseb0rncwYuQ0YlGU30ofZWY96kP91yUF5vPQdsVisNNzfK
ayewHzawfDuGQeQjL/e4H5ZVMSUR0OyLSZt38idm7Z/SoFIH/luY5Js6kl7iwyFEOr2BkFYbKxle
LOB/j+EDxXwZ5VUvdN1dViwLzmrP1FTPO2MKULobYi/SIG3VvVb8yB7++XVIeX6E/a8EnM9m0+Cn
bRWHwHQBOMJ3zFP5JxUs3oA6UJYE+6l1pQ9G1X1nNLBah4U9C0zhTgll9zWxhAqK368m5s85+pIE
oZ0BVkYFlhoRmFiGgN1COlTQQ+ln/Stnfy8MIfXQjXBBifKSer5GNQBxyQhJOfeh4zGqGarOxW/M
0MqjJJIAjjk04CiLFmtLxDs3YuqP7v68w+zLRDv0fEZtng9MIE3G57Y2Kb2vBU9PW8kic7XZZsTg
Cqi+UJrYGyhYoJHNAZ0GErnavTVxX8hMUvL16RNtgKP0n8ehch8RFh9kr5fDQk8PI7FqaFoMdGRF
S/7BFt4nUzNzU40ubkmKCuivaOzT/tp1pcEvzDzAsafekBWAeczO6KnDIfd+9hCW/SqL9kb0As7a
YnbrCkgDGOCI+ju7Prfpzj2HZdtZupOKo193XRLeolr1qOroKQJxuGhy1RM97LHYTLGHH8E6uBhk
RRLmMIx/VKqTOq+wcEa2oo5lN/e92MVL4qTdWWKk/1/NjlsDZqZHtXfb03CsMn9AAKaz2M78sOVx
seE1CkM+5Ko9+uuGXREYryvVbFn+oK4X3+/n0bg8jgQjOQG+U5vEraKCDtzOQC0AC5eqTG7v6dGW
+ojAzd8Az34xUh7vgq47QNahLgA/wYGq2B50WYkoOVkqs8CxeRjKwBet/3nakaKJejm4Q7gnaBiA
qtUbkSrG/t5HOx63QV31myArdNwfDqZuf03kKzAOeNy8RA6rXyYvbaa7JBORDk3XMnYJLFNkCtWR
wEmRrVpcHL/Y8Cqxok2dTmtcD+ramTjXc3svkZogAj7DjDRpolRwSwitsMU7VQeQDO3K4ctBZU/p
9rtOoDImp5y1+fvxj+cRqsWZ7YfAv47eDTpsvttN58Z6zEN+p5fcecZ91v3r97jujwChwf0EvKLv
cS+nIGyHnOoRZfahY1H//XZElghHPnaEwirbFY6GV6DwhuOqs4UILNjQA8454r2qaiw8XWJTgOyO
wvXrlmSaNNQkN9sXbkIlGGESesWOc7oM2OkzrD6Z+tzcsLnCfUajm9+mbRurZ812mtJ03oCFXC8Q
E72T0aKqIaEy+k5KrmHp918V42jZvD2wBvjqjYE6b0SWxeVhF7rGv9HX7yg6KLtgLL23S0/+0tCj
VtWZk7zKXLXpijPU4WimbIrPlWVPzgE/vpTbzQNp+R9Dg1GNRBd6bJ29DiV6x8GIo5eIarqYnNO2
nliBWOV1QKTTUccprV50NtYoGahzRdFVWyBz3pSxlbabrOGk3KDrhDbBtA3wV88lZ9bOdAVzgbyk
bNTMt+/lFb7E4C2lD2xpMKZR6q8z8OXX2PJKKoDgxJoQMprZYi7NCmlRgh6Wy+i0fvo06xXEh9qQ
Mf4wSm1oi/Bwl+OizCW61lomLfH9H1OoAH5TmtbTOjQWmeMdKL0Jl6o/L/yjFpEbuBK2BDkqz/+3
tqX6PpDtD7CjO0lciy+z6ogvBPhXIvJ2y1qo1y2SXXaYxT4XOzgDGoqLQeM4fHYge4TffrzAFF2d
IdN0FOLNXAdDSR53GZT0U0Z2aqRbKnbc0KwwpMrNjovIJrrQpF60JsN0f9u8JrMWpU0u6PKkTZxa
w5Eed7RJ3N+LC4iydO/7RCSwae4LQxj1sZ5FyCiCAuNMHRbakLl0IkJgHhoaRqYhyJRrD7xaGcMR
csYGzss3ev/BPjfh5HCkY3VMmgKjB/8C4yq40S71Rrxk2Z8uxir+uMl4wTHnP28AusWQYeEsTt4L
EIDxv2ZxZur2GnsU0y7VAAMkpvW+fNNdEKCIQgSWM4P2Pf/F6g2zVDiMgMCrzbLjQ8t/9V8OJD3h
GIi5scyq0JAgxpRUBXp6HtjAKuT99FqC/+hBYhIN2X0ZUm7gP6FHPeDfdgQr4DXpieuIZX8uU0Y9
nH1zGwnzVxi5d/N77JwESz21NGCVn+ywfU+eAaHp8sYV6WLnmrLwws09Tf7oSExXZfuluzozk0+l
+5hQ+38/dAi6NZODo2jh3RGD9GtGflhbKoiTB1rV+HQE4ouLgVnGqw7oIbakNdRLe/kKQE+xVVKE
L8j6TU8o43bHbTewp3qx7FdTWDys+K3cAjeTTtyFfaVst+LzNpIvG4rOLnD1vpHZWHOH9CAo1+zz
FxAVA9VIh4Ysm0OvOdGSC+5QxxSDuilHcbp+zMlCui8OkFlD54+Z5mBBHt/IH8Duoy/pBelHHyHm
0mOkncafYAM0FwUqhtMG3sZbGM62YlVouFnpDdOvtQjbtNBMoy6+NzBzw26PHZsKydsQA0kjJlbA
QwZS3F5oMfA0UVUviV46dEtufPSb6OIM5b0nN8KNoOQk135hvwUqmC5lgcrfvaU54nuxGvA8cIsE
i7pzCMxM1MQaHaJP9l9hXBcHZLD1nJo7tEz1AdS1JwphdbsXVBQ6HvUYnwonXsFEQDuMoUi1mnvJ
sfEbzlcweW20fRPLY2Bjy5J67zaWyf68aXB9b5hv7qcn5RiVBD1JZ5fY0X1HEFvhrUUoqLMvajl5
HlLh6p3p4aK5U5JkhME8OCJSwBVWgngMLdC2ENCL1ItgA9W0MOPgSaxnCyEuiOKIAuG6VSgCB/Pc
NZCG2ZqMJJnHbXN4YruqY9LrROkRLp6SVOUzsYfqzCAhwI32mx7tSgsHKbXkswNG4ATX+QjljBv3
6l/yqaD08SaEmdEiCe0UIaRfXhlY9dyqNUbZGT8OmW6czdtz2QxMtOBRlcwP6V0aaysrWMJoQIPY
uv9aQwvgXesIXR7HxgxZ0yND362vCDqGL6HKF+ZEcQ5bYAfPCyu3OhliDXgfHnZANm1npdyC5vie
3mWDucOJr3qLf9QrjDnh+TymuNdHil/3xqwEtAQvGi5zzKVn3voaytL+MzPuvLCCDe1UTJk5QvaV
Kub+dfIz3+pbsai1378zx+aGJiGXou2lqTuYpZxD4lYNO/dX/M/65iLgbqBRtKmiUaOorpq00R4z
PrHCfHslutKF64tTZW5IcHBBmodex3swFUPBrHFjPP44W3KrnXs469MN7RPTzvB0HbXVMBkih6qG
Cp2cnhgoMNZdHq2gmqyNp7K1eJPV5sXw6N/qUQjcNqTfQXXiWFwREOz9xai6g7/ml+fYOfoH16Hc
Sc0m62jX+025bLjLP31qz3E7A5wKyD3d78Rh4ZSt2TEvu/YA66wUdrCxtbYgCZ/Q8Lw2nnmZ76Oz
E0hv4JOK+SXkgLV9yZoWXKTUnS8U4z4Azg4mecY0CWnYcGB1jt9S/rnXV/0mFTRXlueNPu4/7gAw
D9P0L6dJaaA9aXhtFvZYFrgixR3NwoPjYT4fFdkLw95gkxpFMV0EAOdtd6xhqDvwvzwIZSL3w98/
0YvOtVRZPx46Y2IiI3f1iaze9FxuCLlUcK6IZHw5AsuPa+7ySa25fIfFrnrItdBY00uQpvYISEwQ
hu+a8+MVNxcrz/58Cm3SljzaxysCefes0kQrWwxp9+G2mr0J1h9p+getmttj6AjxspU1G1yYRdbB
bXtmN4iNuD6LOoYTUout9te5OTFLezNZO6UCacviQF5NzZ1KP+m1DkBm4gIzzTFlfQvSIVbP/k4S
yPHIPYvP+QczdcS4ITmXc7jrIA2/zV2TOfExJwpwV0thR/UysfqNPazBrQi/vLl8+otoKnCwDmex
POR42CB++pe/1earx5Zict0bqlXg5MNJjQg0hBcLGN6vbUS/drVSclNYwXqzv6+SS+72XwVHGUj8
NcuyHWVm+Tu+SCV92mWuBdisSbyqwbR/PXIkbOasJ06Ol0ySfWrnvZUxHv0hazxNJIa0KrxB1g7T
wVTSw3vtd9DXot+nINqzrJSxK0YkjhJOlUSUFWmw2HV45Mv91tpEMG5lk8HQEoOlkIM00Q9O7QLI
JNX6Z9aIsELrW+ee+QCR6cBQO0uTuL8c4ayMu4vw4mQIR59H1/tD4fwwWtl4fwyO/QLDRq+/qolK
dfdqRWTpu4vLn+xmC18yZZjdxUM5PX+MOnD7Q6c2Sa9TWgORglWT/Kvet6gAyHWe5kbhV4nVGIfI
x7Jitcd4UDDUsbc7sucVZU2gMNjQjXI9O9qlq21CHjy+SkUyinHhCUWokNZZW8Vfg+MSiMxAXzON
/Jd1Nr/6aZwYUlyvZFnlg84CGpxrTU9RBfde/pGvDlWNrXU0Gl964KL2HoOxrqJzCQrkkfBcJ6qG
/z2lB7plANx0IekasEEImJSUIE4ti40zFf++p0RaT+lcEJ0Ej4W2d4PN1/L0lTofXFWxYMMFSb8l
K8cflqbRYt1TECanV4cLbLTAiMOnJaD5qST8u8YPsRkzm/2kXCh8+G2naXAobG/XZqS29v6svBUM
p2EiIBxOM3MgE4L+dBq1APLUkTJRHPcpsYz8CMAObBtvMq25535Prt4Qt/8Pk8SvGczpToBgIfdb
HqaTzb1UuX6bvtCT/aC3R850jlNCYGdlyerUzKviYEntUXn868Jl7qm+BPTNWiGzy6tpGWxV2fZo
nNvsBkIqnJXKC5YSH9LpfqA5cpQtWUeQNopqc1o9qRDCdIN+hXWFp9MyE38WrtL4PfDJcLgK+n8G
lTkACBOBQ8M0PPmI+cA1RdtjXlm3U6iRLbw/KkdtqDJA6iueOm8QbeMz7GlFSmQzhdf0pHAmcRu9
jN1RoqzKiV7z43wkpDeHqYdVmamQHfEAZPJFk28KXDj4cDGtiYyKWF8xX7RfZqy+sAD8oDg/oUDp
ze+PajCiMjLwhIpN+lb1fAGWrCmYMYfAFepZjqdfzEVtzXPwC0v3P7TnLc1Nc250jERIkV85s2+r
Wq3phWFAV/YwtM5x7Vel2nb3PamMohK0jIiRReOS3pVrh//54MD2pPGscZen1Gg/fzEdReWMhp4f
d8LXzB/433KQSLm7HDcRdqtDc/tufO2yv/mSOOasdktHJGhaEdrAYtXL4VsEbAFhluK0u8TgIgQx
wwupbpUz912VKwtfkJif8zCCfuHdorbA9OnZVaMyIucMbKgGn17xZ2Gsh+PYMt6I5Hu4CBko0X/L
4eYSNYXjWuFeiuyP0YThlGDvy2hP9eG+RGBJMtt60RG9MekrURYiVyDMdBxnCswhTHkXiA0lQqQ3
ModGODdqRW42JsxQDOrJZJ1OxHH1i81k0+++NYqskLYmv3jXFuRFI1QVWl6rpios++rPT90yuyZr
e9mxH4VTDw2g1+bXvUp6DqXsYV//iez4ib8ocsXpA5PRHPVZGj8nUee4rLqshNvSmAWFih3oRs2y
tceU9NWaMg5pPQEDYztRnEUltZnVq8P7jEqUNvu13B9AX58Dw46OkASYzj36COuqyeBDdGRHGS+6
kfZlyKECybZp+gaPWByliwWf729xijUC0iPx/C3OwMAQhkSpy07/WUGDB66ENd2aIn4C1Nu2Rqdt
RsdnwVz4R01+vh37fsn/glf4o4T2UdAgyfWfoiDuSU3WkQpuo1hTBFOJGHmDplL57jOj3ptlELYa
RuZPCqzkqTSbZwi9RbQSX/PPVTHrwI8E5ruE7zWT/k2qIpbGJ4kwnOl7ayebV9+2ZcYUB87KFSNK
9cg06LbIoMD5ynaKY7T7Jibc5z7/wBeVTnJOqCe6Hz7Yo5/USzoE8i6pRntn+NhKOGSo3lSd1fQc
4lDjqeOzZsObI2SwJ5Ch6yFuWpGk1syeh71v7bldzxsnj7+OnU/8fTqVt8NVHyFe2m9gFJejdEZf
kjNavUSULOFNoY97yruffGwq2W10k0QSHJuYw6JOnmDbiqGaWs9kbUeGenyCCfnCKqHROQWch15T
0hraPaFL4FoUrth6hWwiAJZlgpKKmU49O/leRQAjWHc7rLeuVRzWAsiv2iQuEcNT8JOYx94EuoS1
cSgpu2aFQoDo5itwybQ1q8B8XEwEfyG0/xEnuk4+oDZmvQ+WaJbun/UeHNJx2PD8tWGILmNB8IxE
Ho/9TApd0NI7emY1eTcGWJcHiZzgiXT/UG6KUtumENIbspyvdZj2KiaRYCELsXzYp7I7mmDhjCSV
4Fuf+K0383+0d5WcpJue7dNfmYZd4uBV6VYgVQ+GQutzXKQzPkfjXiOn+drs5IsTfEwosZz0/yQ4
zFGrM+KDADu06WpwS6cS3TYzXS5PxOVRHGtkBK7Q8uYTZ/FWuYgUVmDdqbpGGW5r606P6DOABC9v
54ddEzfYJXMjCewtQsa7/puL0oycPOAX+TeetjKuGi9djUGt734Ue1h4EyDzPjru/wLmq/eXJbRV
lrhB3Udo2AJoAmDC48tFo2CUI60yGoyz7cPHEEiUx0Zek15ogTr21G8wniU8gQnqACq74VPmKthu
ztOre1+BzqcTmplji9/DTzdFFP+U1c+UvYDyOote4VdC5AD+Zqd08sUpxKnhPD8rgKrzeiWAXBG+
C4FJkvnBmxX6qZGdIWgj/hGNXyqHgB/IJcAFqjCqzhy1yiI9fpvm3909rP9VOLhKCTmVuUEYDUql
D1EkEm8DaykStMDUfOfUoJjuzeLucOxCnSVYd4Uq90fpkvDRumP5MeoPZqAxUebe5Lp+L/u9hNgl
mSOMz/KUm65Gv+MjjPw4v6r681gqc39vjV945ANqae2ZbHQsK8+QRIkSpAxFJsvvRT9n1pJtfRNE
4TXmn3U0qSjFGDRvzZay1PjyfMW/UUyT7ej1KKpRprlhp7fn25SyfpnmE6bZiNo4npp2y4870m3a
mcN76mhB6bAGIXgC8N5cwADb6FZty0IVeOyYqZEJIzq3m/YqVpIoFn4dxNlS/Pl86GAMH1+LkBRC
KdY0kpY9pSUVWrJgZ9EOrlBIZ2cTd6XSUY3Y2CwBJPetuYaM5cN/JIdsrltR/Lw+77qFbwz7ANf6
Da4Y7wD6agBxrCsAjdOsxHP94Y4k0R41o2HaJv+EkKBISAoIWZmH8Qr9REcLPPUFQJx2NvSq3hF8
sumunS2SPsWajo0pC+ylNPdSlHrvcauBaqxV58VpRg0O9t/+hbOWHx9Yzg92hqIxy/P82YTvlAY5
JgZ741kBFG62VS+o4pH1Hubi30t6C6Yd6TNULfIiK4qT4+zV4J73y1MIHaYeUE0Gu7miVMBUszSQ
g9FIjtN1TJWvu1gDYo90h6p7b5SA67pdfqz0ba6RnkjF/Bytr/LSkfEdJgrOKjJaZ8XJRxiQu65X
lUaKbfzMs82u92lv9lnfZoO6yFTzwevRApaOZMENQ2ZW2FgFMJGhes3MOEuPxCjEiX91YcaZu4d6
l6PYBnMDoQMi2BQXrokhgGUVPSHGUEtXhzaZaZyhMp3H+SCebdi+AE/KMhBvMXG+G9tg1wnUUiSO
18uJllOs7DbsVgKUOvjWnv+qmvNtSQYD61Xm4zfe73xVAJ4Rf5iqflqje6PSEmolWsGCF86Exy77
oKWJoT/YMLFOSNFqOM5K9bJfCceeP1mbOzESbVrka9HG75THC1oD6FmUJ03fBPwbxDfx5ssEHH0y
bB3PHZhlOVGbLn0tesOWTtXpp5W7tTwLWOXT6UW6UDcYwPFUfH0PsMI2DtQKyb/fWYq1Yu8bhiG9
qMkV7hFTSWHiLlwt/7j6mYL9vNV+mFFJDfWEHQeTtndN+3bi4xmqyf4IuLDrOIYSlKpL4/YyBH31
7Bq1asUp5mlUY181bzcpteDk8tIB/jvrEWSqBp3aZK18bmZfggysYK6bWPUT6tGu3O6NHo09oRg1
6OsaAEHh8F8VfKFc5jdC/zTEj+QsqcrHcjvhAX2nZMxcDUgxAYLXffuXCIFTkXuq3sGscvpBFOif
bZWLNJp2K6IyJaZpBc4YDm8lfBc4u5dWl08edEWCQfYkIXDqL3X0qm/YCn5NsrLJdo/9jqWAxvTH
E3qOgekAzPy9hF1HvIQYPwGkb1mlaUN2oYaYQB8FtOXR8QtNqK0FRtiqiTshSTfJ6SxIZ4lSCd//
PKgOSGY5CDHwi8wrro+avMZgFM0eBMHmDCv5+0v90se0hIJMg3dboKFOh73dVAqmBHnEh+mWdg/M
AgsG+u76xkX6w7stG2fTpNngLVbrBeAb0MlslpkG32li5qlA4W7etIx1v3fvQJ7AzsSk9zeBqbwv
nVgd6W5OrU39pqx5Ae4Pu83qFqZrTGXJOn2r4vjILGSqXOpKu5CZcIfpGXkGhMJYvx0jQ3cH1RVk
YFtOViyLOn2IyCvkLlevFUvupWOonutm27xnRe1HrjwEwb4D/b6Bmo5FKLWcDm7KRzfXRgr2Rdgg
Scd5aeknQ7Cg3vH6nZm7R3y3FIiQAQx9VARP1fqXKLSnM0ky+uDtaoccZTWrQfijcVKO1bLCnucq
jOAfKgkVVcl5cW6DqdyHatwvNRxlG6kDfQvVL9HCtEiEWFzLnHipQRt+a6c9HOyhNVvUHUw794+G
WZKIacd6/O+wCEqTGBmZ2fUdlenmBLO5BZa7Ik7RnFKvOYM1wFUPRWP2MNiNrB6s2HfU8WKrHqgg
bU4gJmJzZpl20QCfDLaKVwp3x5c+YgY+TgvEbLIO6ZZNkUJMOfv18ySfe7gJqle0JTVtBtsfjCLE
I2bM3BnMdTmHUneMU5cUUoA96xmU8JSHgcEQgzXgH+YDf0sg5P1NOovOCYwR+pw9pL0fRQXvNnee
2Znpt+9wr0J1LT4knNCMEweucYx++g/aXLeumzZk4bLGLyNtcLy6DUgQ4s4emEThDwTPMJFFxmki
GBLDR/IGpVP+k/7P0lcX1IydPu7XeK2yVPurogu823hq8dYEVfLx2flBoN7l4+7ax/w/tFLLmx+C
7d2LvcAfXQgFdt+pk3h/PbQvwqh0HIUIagdxZdySOZwj7N8GKoScEvXtWwydwahK22l07UCU00+W
8q3HgpCprXIHoAjs5CU4I8uS6XXDYA1Y9RRCYRXMHPZTJvbza1J0NfBRKKXz7ucjo+TbTeh2ZWre
GkKqb8XJqfQzZGBZK5yjE+a90Ko3lInyOaDDnKB4S3oXqYlaUPIbCA2l6jZh4GBgKDKM0LVlhQZ1
8StesimvFLB5t8LhBVL02V23gnbmOHksHLrQgE+utEHv6ZD6MkIiKyFE3pmf8yJ/BdqHCQft7XNa
OVZMrMWWASfj55m2vBYkkLcoRUNKj1ohXW9uAnzihuIuZdUIEwUxFLCZJTit3KwCL9DleYvAbW06
0Rpa4D+DxGYJSZlHs3y+tWkUGeuqf3is5RUFOu92z8zT7EMyLw47q6vMa+jxxSQ6azaB/SZI/UX7
spTgIUHa+ixIR/ADwxLSeCPgJoP4RrJnwqvzwq+jNR6/OQJPcIYglHzHJeYwNA4dB8ZI8B/u63mJ
34woa/k4+0oBthO8dEWGoKc6eEkBUT85NIfW/sbyCMJkQA6lNh0ba+ISIC5EFcEF5t5/CFi8zzXE
T75G7T9BToINcm/VY6Q3c2CbPIAKQj/5BwWM3HttS4+Bernv8xCE1RgOLxChla/lsIWXIKNnKBfB
g5ObQScmsKE7jOfI/Uy37MYyvjYozXvzxe05/9Gwu7LwjLv0PHP1x/6wZrZEGi79TWafmtWEY5+V
yk78+UA+6gudl7Zh2WpGDuqdw5eM8ZtKpVmcR3vKRg3u9akuo+XUCKmowuxFf55n27fTqiNJDOnl
/BTlzNRdGvgyeexI2r4U1ZSlKkipzEU75SOWE00bl3cb5ur8nfiXF9yPlmQLRH8fWipL5i/E8Wi2
DhupwwQg6vbfsVrNFKvLMy1FQh1Ph52ObNEeS62BkewFXv4O2QKOO5zxmuB5O/JTu+LzQUSaTa/6
QCdUh1bLAqYMcWKbr6/nJn+mTrV2oECmJuRri53r2v/Xaz6ic3Fz8qi4jhy9E4jPd1YihfgsrKyi
8G/cMsbk/VAXdhj8eYNq2ian0eo+lfozOpFbxg62GQHhvs4XPAzqwQe6TbFA/5rvgwQ5b4mb0SWg
MMMLWEZT1BuTg02pyXWxkF06sEPEYhWhlDSgYZG61WQ4avutrLCW0WQzMtD72WJlGosuIFFtNMg8
tPA2XIin2hINldRjCMyFbByz3vfNXTfCKDGUhw+YMD2ewnG1S8YqxtfjTprl0lSs0JPiuAP4OG3r
KXq4bWdq23x8f2dn2gNVdADhOxZz3rh1Ht2dT4HvdRtooYYFXGqksK3sHJl7462lCmXBfGVN2c25
4DGcdww5q3ea5EP97JMYXL+fF7VdHrI+ggoA312hIE4Rj2Piiys8Gin+9i8rHwGDHNN3EJcMgc9k
MnEUvUpj9eZyzHmoLxo11yJgjamji2kuKm49fXEKylD9M/QjNyqLv9n/XaoTLYOKSlWyVHJLogdC
ouMUOXexKMwRLbmhowtMMQGwTep+wVIpbOnrZ5bwHw4c54ejgsKfjSU7+8e6Q4qNNhNf90fvUC/2
M2dOuZtk2bzm+9IRWWnyjJeydXBL3Y02E+NZiqi8HXhgHm99KQy9xyv32ZKIVdFbx6LCa7svu4eo
lfWA7YYGlIuCZDpcDGrOc288Acuu4IRzV94+5GoVSsnsODZa9iowuo96hYQEp84NAdTg82egAQuA
K2mmOvYFQFbmD2+boZlA+HT+xcLvPfqttpHWD/Y8fbJxikpqWC7KlHWXRrMIo/ggdHe9NWVlhxfk
0T2XXWw5xBIWaK7d3Zd4+7b8C8/DwCWPI3FpseypITNlnekTq/GwY0vNv2PEKS7au13Z+Bc5B62F
bDt4Rig9tkKsvSz2eQOmE4naEgTlqVxdoFbtG70NUHT5A6YX0zs6YJk9MRb7mVH6CS8zmVuJyzVE
T9nVZ2mfi9DvBGvntNjAQGFa/DPcVaOHy3vOjJ01CiHGnQPVhTSm/3qA1D0iFo3ePcCxLI0cXJBn
XHeZDus5Lc32w8wzwwdzFe3qf/AyJ5PSW2jFpc6dl4t1nsH7QuYq+H3QmrZ/ufSu9J7apipbWlWL
NwaFzzyd2Zs9yu4ZRlXpd+sQ40FjxI222jQcVsnU88xzjS0qJ4UzpE6my50DjNXNZm22egW+Vum0
vCHLs/ciDkKeiLEnh7vCD+nGDc5ztVWaLZxmEQGXXzVIhR6ttiq8Bhc4u/EOednD8BaWPWJd1P+K
edcTX/C0R+VhyZL3UjTGGNx4BzeMDa1rtF7XsyzfASG5ByJQS5LMj+6tyWBqWwWNDaeVnD3/4ZHV
YEglYP0+WEebd7pj3uwbvhukSOxe+liZlMHpeVcqPdiTKOhFWItdEXPikQMF+/+20HHRw3EwlrbH
u/jvPHLx7xFyP+NN4pc3xzSRo5T6K1krNEb4I1WPqSqabvBuB5wSvhJMRSLMG7HQ/26QeTJyo+Yw
RmG5dQEOog2oAdlRdQDvx3zkcgeMF4tbWMLA2O2PIACftoMcgx6JPmfgu1c93z8Y15k0WipAr+u2
my91jA6AAc+Zpn4JUamFAcF7iekFWTdJbgRr4aSaaiXNXuvnbghhpnuJ/H4RvauSiqa8MX7r0ZAX
b2YSLBqvV7+GIgDZyqeaGGIeMH/VQc3QMLkomJR17qhHstSCD0UaXFC80NyDTJMHXKsmFgtIk3wd
M3GX+B/GEFx2FuTsZSidglUgm/SxajukYEXBFKkum4Umk1CTnEFbr2NOOvo9k17UDhq2nMjNzaVF
KrAyP93VzCf1xiQRAzQ0UwtXljCvq/r0QLfZvSscDEzQCwkvLcDTTe0VRyd6qXLjE84c4Q8+ngk2
t4CMKkDicGGevJ6xBMV8PHPXT/L52978+K7nMYDXRYFh/sM9jhx+aq8cFDEfYVzvWGzn6Vt+jNVc
WVyf3kR9hyMSRAW/NGOmyqMbRySYuOctkz5oZr4sktUSXS4hlh9BOiXCaugkx/NX4bAx3q5aeNE4
M5OdipPhqudq/JPM9pVLPGcFR4R3vIM9gCntnXOe4ARuwZcX2v8w8Jd8qAcJpvKEUQPEcn7Yw1AH
R7wPD+nKzai4z80SJ5gi+TQqagTotciAxZ7z0Qunxf/LXA1hxuVjpTXIA6V85lNGYuY0tm2TLQZR
9SdJPMkA+goTWqOGxLLAiRWXXIyGrvj5g9acvYtr/Er6m94IBuSPwHqTDXKNmw5u5Eh7Y89ja7fL
XoJexxU7oL9ck0UGypfACKIVpglBtPmTZ27HoYZfG9+bPfPndBPaQke9B/GkfJ96ncZVzIJEiWX9
xL5BAV3zXpvfHOq2WnwbFJgwfLsvkbOC8JCdHqF6VGlohC4Lidj2lowQxD35dBlXskHcKU7PO1mk
BEuFsohHFyHrBamQytqD769KQGB29vgkmvwIIsyCzFsc0Qv7I+/a6bMY63uV5FixD3VyUnU3a6t+
3FKClzweBArfyWUUPVn2J3Rl6iYyW2J804KZR0ZyK1TQdjV0GsC+g0waAAkx/gQp6WEs+dtUq+Pw
w9kLySJISyS/NuRyLGYw9D9QBqYsvGDCmuBjBMyVmAit4jJ6t8nJWE0n0WxISlR3bmA1bJQ39L96
ab1C6nIM7kJeOqsHrlvMKwlQrmzCVVp8k2v5b6Km5FYhpMRwD0+ZTlwO/7Uc0FEWx51Cd3zw6m9x
4LeNjdQr2YzzQIZ2fivOGQwp85NPdzQN7yOFaUWlSl6FdtWHjlyDEIKJJi78iYQJFosH9X7WbI1u
egNM7HqFfoKyucnEulZ511wR3tXlIIPIL7m0oC3+X7otHnqYztPPqCfApyRsZzFkmhI5fKh9piGn
8Ylwz5NmF4llLm+zBHoWdRnrHoVt1oMbRwIVL8o2EIYXxs4jIjsbN3ZhwHmXCPb6COwGS3l7Nuo0
wUZS8CptIQblWXoKyyA5MaBmKgiakZKxqUF0VnSrExjtdQ5BGc51D6Pb5h6iXZ95Luyyj5qUix4s
5z7ICTDGE+2SlXmjh2q8RA9F0MUnLOWdlNroAK2JS2hO9w4DoHKB/WIfyiN6+FQDfeRlmnVXHDil
VxM6R655b4r5R8zvqMBB406dDtJ3WiVn8yj64fWV237mM2KJUa+vMYusaJzVvhHDxzvfHDxURGUa
uyiSO3ThxTUllwaHN/nIb9F67pyUaIXFxiB92xy+nQjbfpHLcgq3BTTHtvSRvtK5quwbL6JHbWHE
0nDqLO2V2A8PGTl+5VfspHHbSTgLI1yXjGEebdIHBbTmXWm7LzfnyKlmdam8Y7u9sNakuBfx0/id
hAmhn8zESHy+dDUsixbjHdoR1AwUZuvuxViDxBiiP2NKkUfwwj8fVSWiLz8gjnpazoomKegwO9pD
iUctnZcQCxfq8Sd/NG/Ysjv2ghiluIkKIvyAhPOX0M94T1ggG2GUVJ+w7G4r20ulJiCfiKh89yGp
DEDD+LLwly95RehiyGxWmSzf9Av7Il08cVx6ZaJa82OVhwxkDsGe4qb70oVdXSdigF404obRnV9s
8C/Tto4F5mxGHajXurJ4ySE5O+JIXp6UCFeakxndPNBDwYcZNNHROcKFgu3zVVYQZB5dPodn4ctC
RJtwxOZED4XYeKoq7RqL2YLPtlR2go3CNmwPf4xA8d9mUP03oOUc8Z3DCfpZ6yF6pNp9pjEXpabS
JIrTHRX15wlKWkAVQGDC//HH4UE+ZnWNqwXsJ3dYsq4N49l+PiH0Y45eO0E6CT3QxIgKcbwBmk8X
Unaa3r/qano79nrF3NaJeNJYA1R0Hwn02qx+XdpIJKDBeZArrLDrqlh7R0OhfrJ+DJ40DowF0qZK
E3fkDKpxyIgVPTLF4YkEX62Jsu8XcXj8Y/vSD5T7Hte/zOBfywX5+7TtEKIAp7bwz5slcnZw1aD5
DFz4tmIPK03NpkEpA2o5jakiJsn9KrzPxAYPiPhfxKn5wkhTDGe4KU6jC0Q29q4u6LyeQtRM0vr8
x7hbDY7GjVFQP94eqmwO0TdB95PM8zamfDLRWJmac6/5kVPY03NNxRWRXJGXP8vLSWWq4pN6o4DN
Y3mPAhf5hxK2oR0XWoAffj8VIoRbH3GOpYLORl1iix2bo7bziofzCzwz/x9riTCKByrEmGiL4fHs
AN8n+8wDjUex0Yu59KOzuwWh9MbWh2QHN1nPHPI8S42Voj3FPH3J0R/vediPGm4yD/JvsuUufLIl
embVorxkSFWDPJRcvct0mFgmfzVhW8TW5Mbe3EtLvLZ3Vakv461unDpwa88crLHdgmTD5Etn1Him
2G68al7TBFRNJNghzsjJN1WjQbduYCOy5eJSMl46WHRPc4Ht2/0jxBiuAUAsK0rdROx1vzkHBBBe
tJt6BsXJLp4C9W8qNVFKW6VNfY9uQ25C2nmalWngVK21FO/b6zfqCqiXYt42Sw5tokxtIGgcmz1Z
irx02VRN0QoSbfPh+39Rm6g1u5CjsgvIakpUEPwYrhKUy1H+TDlpbRbczLrHHQXujwPyflATtP2V
k5D/naZsmyzlVA5lzQdRuw0Ej9vNv7P0vDor358u4JJ29fFcPY84eAQEK+syGFg2RSZ9WU7VIjy3
vWZylBlBavDMrnxUD2kwc/arXfyB/RxsghNNUQTLxo9/ocLkPfGx7Dsac1d2v90a7ajj8586IO6B
P3kUUkj9j0H/dVYltKDkacUwJtNcf5y9EFAmlqOGrRrZKGoENuKId4wmnf9XgSVEm0mWzGh43Byi
aqlv2XEYp+zKuKUxuQL5/He1q6cTIiCm7QjI7wEpFT3Odg5eRk0cqP86shBEn0XlOL0DL7mj3Ap+
637Af9wJZY73rXCR6gnR0oqOA+P/R0wdz7SIUbpbbv8uduAvGNBsfMgtc70+0e3VN12EBIJvf7Od
vtdxc0V/P4NEBW/Y2UqE9ukIRurCX4xk98fWYXnqvT3WQYXwiH9pEpE90QwDtkfaSCmVtn78kCLy
bkYJ6GdSK08P41jh+i5yXvJAuyjT+gxeW0MHrwBTZWCzEGkrWJwj6CuZlVk0q/3+/cALotzzqUoz
ih/igxgi6QJi8pTvRn1XWR/TA7bAOIVaCmfgQhoRuxhvCkFavVxgn+r+jnBlptqCG/xguBS3fml0
h86dROhKkYdGbLqrDOcq58BDiWNeftYPGpDlv/mUMC4nSgp9+OAOGym5Giy0rXXjVaYuGaRN1a4o
HLbtwc+ffehHR+KAJZcevwUtxnoORvC12R420y/UvYz331vTOyZ2rIrmzfv7GRz1HuQ+vLuCamex
JShGNVijB09nphHN77utQ17OUSydd/VzqQH7/k6fMYrhf4xnj7riIoaqPZ2qEDuuiNNrZrrVwfAt
nwv6ebxDOOlCxPO6tQSwAHtu47B4QxDaZJMQXL/j3utCpehdFhSapKGT/iPS2PUtd7FKIM6dCoUY
HKUABe7l6/TkAnMm2Rmusg8IypRifEjD7Nui/ez5TYHLeqFaEnu3Jtp5yOGgveH9AwUPk0TW1tK6
uzb9HK7B0XRl4lnbbZVT3eU+9MjKo6mZVcbB0s2iDVPgpMw4Ap6hQVGI6Ye4kdCv0sGPxt3u9DwT
yLcKSYjd1UlIqSmmKUxmRJYgf/6BvkSRm9iJsmR3dUbSxhr86KFnm1cZkfTXRuMOEJJ7CxJj/8Dx
kz6wTXUNqnJck+yok4FM+nDojLHuJTtaVsyzwTaVOddcyQQoKriMKiA8oGoKM5too1Yk+6dcOGGg
gnxR6ysWixfqicsZufVe3L5lna95rbENPsVH1QnpyxpkDQiFGnVyFpZxB/RcEJJm7Jo5gScSnoo6
B+xqcV6n2xBprx4siTA6CJHH1x6hxAvncjhZ7uSliZIdTNOtr0YcagRkRSlcgY4aZJkoRSIR/QD5
YpCd3CLWcaFnNJk+qYL5W5AYb440f42tzW7yseJ7zNNNwcrUzvW+2ArdmiCFAa8RqjWBwwlKx7rg
/oxQDJgROQyCKNf1HqlEqSOFtWSOCZaahO0GhJzDpI2hRnwmrm8LRmYnot4/XWxJza1qjE1HYvF7
s5sF/mrMDvjevdaY6E0OwYrTT5Nur2cGLx6vmHFIuRpZWQaWQH88FsdakFiQixLXEIcugMX3TKfh
cFun0VpKZ/qUwK8DW6TkjJXlwQIVHKW2mUk1pnqsgC8PgHuSEttGOpR3IBlO+eCpi734u7DngDUt
c2W8Ce16LZ3ZIgZ2e0TBM54Vhgp1DteACNEVGr+DRJTKQqD3lxsepXhlo1nymiSyXhsdapO+A+Q+
5ttQf47eTci4/IHTXrHGZP00IO4k5pRGLUo3Hw5fy6FkFskuBNkDEdgA8G5nkQJw6AlGM3WOPOwR
jbmdnpyiEUU6b2E13NGQUlOkDeJk2Ki4qX0eYbKRZxEsi7Rgfljr4sPghx/5N9Pg25+pq2ThTgSU
88jxBVdVDqe1oQkdHRByBprhFhg8JT67TjEw3X/NGkFJcFrDsJfkleBoehlhW1ZGM3GqhuXwnzs3
1jFqyrI4GKbd3kL4EGCdQ98nfKJdaatoTCv49y2kAWZGRb6QEREJFOTKqo636K+sXkjdv2m23AJK
SlS+k63T7cSwKyHcDVbJpZvpGRt+/tGb9B4qSmpNKenL4jpM6LJOocN1dvOPXkbchJNStKimrXhM
3C6M/kVfNKIBLpCeafG1Qz61H4WzE+vpHKVLqk+VSJYzSlqW0T9rhJdjKMTFyVUMl91RBZoVv19U
hAKkBweI5MVGPJ0KollSGRu/JjRC42GziHL9mAtltLpPk+dWlQiILIXzGyuf1JqtuGQS4mjA2meK
WvFGU7gVn25gs3nk1a7HtM2MNGoN06pzq0E0zeuhnpy/gOORe8p4pwIdj8BTrwK8DEJBiZL7mBqH
hmyVxWR/YaanC0qHuKGFwKvkjWG6LfOsckB3YwcLCRfTldH2pWbaUafQuZTrGqysZEsRK3NQaTG4
24kjH33V6U81qNlugjWN48zq/Zz4zOX0YIMgyWeC1+WIvIRB9AJ3RVvnFTzXDUC4rPpttK/a7jda
byEn8kesRXMabVGUAQbfpgIaCdhhb/LByu6V0AxYSy2unMDNZLHiBaQQn1UsD/9UDDm7uAe12/c3
l8A7Api/InPqmmbV33Lb3bc6kBXaDyl8HD38xicm9ViT+HpdA3QJPrRKzNe5v7jQEQc2gexHtGw5
BFcsjFwJxReCuXfJK7rHmP3qlF2Pc3kIBhxQMJwI2X4XKF7tjPVTpB56Zd/G2CyRiDuqYy593gnU
ujwUX4RHN1bWwVWcjCj3Y+r3OwFs+VAT5ubxNvDX45hRptIHuCKkyu2mMtWIGVCukZTFVPyf+Xds
y47YHcbuW+DPxGNLQkrzuE3zXPYrCXobY/8A+DbyHQ3uZBJxGxthfLzeOJX6LdzAp56+sCBNSYIV
JA6sMcSUulOUrrET6D3TvB4s9sXjLOy7UKDiL6FPS5ITuYovRSlB9WQLa9xNoHG/f1MLmAuEY1tQ
0Ru7bEF7nWfgbQ892g1J6prnc7oCsEWOCK/2qcaIYKFuZmWqutKMwTOQECWKQmvAWdS2nQRQP9QI
iYjyEexy5/pjg1XS4oT9OAiGHaH9IS/QPqdX637H/Lywt5sJoP0UzS3XYu5U0HL1kyCPwtxO8Umt
h/60lVo9ZvlQOSE/rekEup3XxMCJmca3gFfn0Pqli755gq+pwt3PN/UTUszxDesXq2fL7Uaz4X1A
f5VtgXP4ogYGltVf2zI7IOhymi3Iq4FiOp6QwSxZ/UuUmFRg2GrB9dHuEJ6UzLFw2PCAI5E+pECK
rcPzt2SCPgdbziVxISZyEXKUdw6O6xndggatR2zSi0r+pokIDr5YQYAyaqBjSa8QH7tWKqmgbObi
YEBd0G1dd2QvTXI2fa7YgInUpIM91B/CZJ9u1yxCjaTLrUR6Wg7wwC4eglLomslGdcSLdSRJ+P64
XJ2wLWfUDylaIbSkqkKS2QnfJ6MAV9vlE3oASjKpM3NeXH8PI/njYi/ok56DrY2A/lawloSz3mJV
Riehk2d2zGZQ/1mcTUv2EuHA8KD/HfclhRspKCN6hHY9ExrSVlo5QupwTAN3iVh+AYzfmJcqAUb8
Pnm/u+LygFZEigux6vWK8/Zf+UfDKXshpGZtfXx/fTSaKrbVhL/Sw5NQe1YezpyPCP7FnGGCbdhL
hBCrytm446XcvHstpLdemysEE/ZlSEm1f4vxmAmXPKQWo6cOruHszPzBbQ+RaZ18aUrv1zL3jDkc
YZ/5gg1Zd8UpLTwZYR8qH94hZh1j/4UT+wD4uWuuUhEKdHtZbAwjxn3led/v9iq8VKhA9ZlM4pRT
c5Qc4Ap9kBqU3jR2TdAeACEAJAoh3ywBss9GGoNoyypSeY42SHOTcrbIxTCTbi6PaDyhZBHlVaRK
V6nM/VYxMA1zv+Sy7T8NEif4HGojHzzIwoPjIu0yJ0ALWYu3egKCpTp/MUBDUNmXHBfTKv69ubjd
TpCsPdWCSkIZhz/UNUlF/+Rb33amRCPhi5LuzG4y1nttU6Fnz0k3edE5FovIzihAMu7BxQ3aPV67
Tlwbs9GodheaVl+t7mqSSL7T09CkJRaeGd9t8jefVN8ItP/vClfhaCjOKxlvmx4x6LqRVE/KBgkD
Dezqh5y/Yz2KyPXTtz4fGNFKqy9Dua7VXcC1XHN0ieuw5/kw4LpaJ4a3Tav1OYEvNCd8BljjYIs9
WaAWbcURyFK+PCwLLki/er75TFLa2icRRIlS4VNnTMgpSmiyNT1CB+KzCQrgyTKljff2NZcCw0Ih
iyJDZ5vpYA9rK0WNpgds/S4gIYTCUbgVhwhHeHKeZAHQt+mobgdTt2fUGd8UpLES4aDTyV2ETT6n
q2LnN3bSXk0gwPfO3wuka75Vz9m2dEo+qFGzvKHmH3nUGjQHgiNw67XerRBEJBo00wOimd6Acgk/
IsUP7hkyA5AEtmRjpModdSfSg2TyKgpxkPw6dpBVpSjS2FYYOgUYpqnvfj8pQ7+sWgMHJwOtt3gr
s1fEoigZl+nTxcm5uF/Xv5xxjICEep/YhsXWu18q0cUjAVWaTzKxEZckZYlZsEKiJczKzY9kwjvT
lbxanhm8KcdOTVtAvMPozBWDjfhEts1J1G4DIFEVG+PE157KSU9oElsNK0PlPIFfOaDlJ0YrcyqS
yz63vidzdgxs3y95O0Rc5TA+/5TGbBXk0Qgxkw0YvJVBXKLu1W+fSpqsLQZ09uqNh5fmvYhfq2qM
99Mz+UDr6VNOlrAyf/bsoEQVjjmrVvJwyGIp2HNGaRBALmxVsQ/k1HaCnjU4/YY8l1zyv3sM3wOL
uSsJT60SMfLuQQxiU7fs2FU672u2F6Hk86paAg1YFQCNFuhUpAM0e8wqELpWoriQ62j+OSdzJSXD
uq+5qnu1w6FEEZUi9fgG29Q7MIbBBs2yn3cKBG7EoMbVZfW6kJMAN5xj2oWrj3EbSKMtqa/z+fgg
+5T2XB6xLPMRTOqOuwsEojaPbn2oCC0tnZUOpDUPNCArw3dT0AFYIgnLlLTEo1I89KB0yoqVHRCm
q16fTiMzo97zoGZBaTinP1k92teTYOPk3SHweDlxgepmloyHxoDm7sZiOLPQH8rYYfeja6MReM+D
Yo18eZ3VTb4pUI5kQODOBhayE6MP2cORo4UeBfzD0IXHsuT5Jrq3z8eWqQJ7KOltxNqx5LHkzPQV
200HxoixJ+m91K9BQTuU2CJJtnXg3G0AgvO6Vg9VUnHfsWxTfnZIPb2qsQiiZT3/vZwzjUlz8PUb
bqUIz0cLlgZSljcWsqXewiVNY87tmxJrn78bQBLry35w+nNSRr98smuo8qy+9T8QDoglWaG6CfCc
gK9XP51sB1oOpHPdwTyXCUuZk8YP2WO0dm5JpVel6XoOnl1EXl0kc1d89YHBHWtrsxoE3H+v97HS
j+66MQPMhkoGIkzzL/5gk6Yu8pUkAXSZYHnzQEvNf/UzimOp80ZjUs4wbvkHhh86BKKniWoKmYCp
ucwgt68bMGkgpqrKR3+9Ir9+LhbIkORjSuh/7Egp2+7ahJQTLXgYXIYiAi9ThJGKKFnONrQvGeJ8
bRTwVaI1JOSrEEAcoTuNmKcrPpf02sEHVh5PrhUFHazEJZ5n7uIPyqad9L+oZ/y5YEXJuj4BfME7
rtTdNYXQ284YWhqLrz80cMXLZBhm/GOjbq6EuhXghdKgKKFPbMeuBXyvzCoupX1Ui1/PIzIGZmgP
9i2lfSB1ZVkrOEsLhJeFr7S8GwR7YlLwm0bSXCcgUqtubfi3O3dR/rIVNL507p5t/8PmcqsD4jBo
x30caVl3gTkAdZJj+tP0W7ILYxH6ZdbSOsWI5InvfCCivgBrlhFnE5/YlfHxfsLMFYSUdMCNeDBW
CiikQYTPkY3G76Lo1l5gIUk5tAGxK4R4IEwRutv6bXEZPgqP4rT/3fXK9zmcIBn3tP90N4/j/o8c
eRehFalvJ/LcrDNrw7G67ukhZIiz7SRkLO5yDD3ddbWVMhG3GXoA9zo2aQtqAj6HcP+Gdo9ohF0N
miWeBPfyeJ5af+xEX5sfedNvUBbVJM78Pg4laQmSkpK0pRww8tVQeVeURjeead5kwhCt/oHf7PV1
j9mmzOMLuXhtfSY5p7T/22OFoan6P0LIgZZ6x4STFzt9QKG65mRQHRjK8CZxp2SfoSPls/rJLs3O
aFaUD1CFyBIKidVpN4gSW7azcf89NkVUW8hPivInHK/ahLaOGdbBq/TKl1eYubfQ8RcLZRqsV3Bs
//Y1u99iJsvJ8mzkY+haNvNwaQRm6xA7SMZlnHQZHV+DiTSfJO70uIeG3Qr6uqpiR8ozvFCHfDdq
EabGhgPNJu4GrciD2LvWVzXYyyn1fEF4zMfNsivp0oBtmi49kpj2nT5WBjGMliBlOOMb2sEzCw7Q
niANSJOTx8Y2Z7yzVTRAGPSUfvpte25akllRcB7+2v1rHuR/XKfNgfD/eFgfQ3lt/LzxZUWFDuxG
RBT9FHpW92bPDw2oz6z+B3KJiGi+Mztlza2i31z6H8v7sU6bcPDNl/oEmymwqeIiadp8D5HrfZH8
fUp6FOtTdMoubA8zrT59iDrKO93ORL3WHWauxWkiSCD/pCP4L9rsDZ68B7CSv0LrAQVnY43cepSi
hPt1uJOeaLCyH95sC2Wc7TvFLKzcaT+ZFTNdERhSuvoBjP4r24BSPig+Q8xXGs29DALFMJuCyMb2
HJdKlA1q+1IiY2a9TcMWmARiLoOt4yIltdk/zIHsaZQolH+/GmvWya1cDEq7TRVtBc67uy74JsIj
4K3lQIpV4YjXg7MFn/XJfb2yhLIoUwW6URVC7y/nibkNEdO/vqYoASyqyXk+LDi/cgFW+ZZX6Lem
qr7tYNANYvQFR6f7VM506luFQJRZR5YNKZ2jhDqHv57H9fq4euTdMnbrUmnJdIG3gFGmNLEzSUob
id+QA1mNF6A9voH2gKTJYrhTnW7lMgM34h2OChTMG+AyyxlYIziX8kl6DM6eV7ZsA4ANgBWs+9b/
cWmL0Qg0Yo8q2i1CSluxX8Pn2BoPeCbjfRRQUu0vPu6uzIZxY4m1DXIBH2CLWZyyKPeCb+6+7JH/
Q9yL4Cph3Cn5XM/Kz6VFMCuYU56i9LurWcUNpbBOiqcaJEJ2ae6tgiwjtaNhasZGuL00dn3DdEpb
yjKUf0bFtyV4Y6+J7Y00OBV9YT+24f7JVpY2DweC8ZmxLadT2jQTKKoNoZDi1VaRRWCbXKVeuhSn
WqzMhZiIiTBWfQr+7ci+AHx9PxO+RanlJY3lqtod6HAWSMXlltF6jDjDnaUZ3jj3JpQWOAhftcNy
E5DnQxOZmdwrlx+utI7mEtRpKAP1JIlLBKwsKnckKRNTUqTYIIkbS9QEctx+hWRvt/6ss8/SGnJo
gLzbGqAtPAKprclyw0tVyT2QtjA+GuHC2gv2mfXvPC9KDdRtM64IN37viERvAy38TNZ6Sefjh/3x
DKVAfjMFsdn2AC3srca1yJ79eYU/IJR2Jzq3G0qqN6QVgYXsgzDlnGyaqL3p1+NY2/6A1PlU5Giq
E8kMCLUD0KqQiWsN8fwOBLEn0DNHhUP4v/9s6pofo5F8Cpf98oR3JtwX2TxEu+tBiaTWnkppohSj
x0GisfwzR5AznxM3b+koGJLZVVMwCSpacYFmgxF5mM9E96cyuLd1bqUPIisVEjEXGQRfAKIo3aBs
lntlmtLx1zT29Kx0o6normsAbTrQgiVuzHR15wqZcfK8UKeg5YB4GXzT1kMLoXByxYfapmc8vNGy
bIN1JVW5rYBBZY05/vs79JT3qjbcdEojOBbYk3bhsVNdjAbajdXxdjiJe5QbK3OFirIsjxQgrDt+
kIhY6eQ0bjCZv2weETU2QGlUSSakCEu/0sVgDP8FpJiNbdKghbDsfqHjvyIoEMv678v1fMeMlba5
0bOY1+lR2wIw+1WgBrd1kfUfm0H845I8zyoemkifDs/015lcfRFD+ddC3lFApyRfChoHHUnW/TR1
SL5VLM2kZpRwNfgBUuISO1VsQ4Gma4W1yxqeF1LB5dvylRdAUJb82Bfk5UAuvxiV8K6XOztl7m7m
e+0ytWbcrKR2hY7q+7v6ciAJodBT/U9EdBmQDPAZI1OVbV8QjUZ95dc+fGJW4ytFIELM2aSZVij0
Z3KbyLertbUed/f04rMPzhTGtC31dKr40j155PDTrWK1gs+TUp6d9XDDVKrAuAwrnAbAOeC/6pNc
NQsPE1vluZc35YlYqnJ2sxoBcbvFY++JkBpah6K4vAR9EWynAhF0XRdTh5bBlWG85W1DjcpXhKJt
iqcuFCww51IgH3+fErQdH/Msnt2j10CfsXO0cs5GkMtxAh3dEPmYGH1oqoCbZV4GRrvep7kLCQaS
62W5Pad4LuzgL7rq0FwViOwCIdt2MismjQ6tYsjRXdS+0DRlurbldm1GcndbYCS6ONYiLQ5CnD3r
EHwb7Fqttwo5kgzZR2mGRVwp996YeMbcFKqpl+KP5pUvCU7MVmxT6iXgGqh1BzFgG4V188Pn5j+E
gMI/+TTKCRBalbU1IAmjce+0qSHAzjxUxkEr6NWIRUAb9hZ0ztTBBbKli/eClrWPf1/jz9d4zPqE
UukD5togPy/BItwxWf34G2kIN0Fvjv52orb4LfG+nMCXLk3j29ivDAomUFkWmIBN+UblOltpAcA3
STStgIIO5EtJ+jd53ewYwwdlmDQIjeeiucufcroBIM/W3snBUUldLHVeMLaTvxcr98Uop3UNM3Hi
aVQ+XkUrv0FBKF8f8SY6MsbjMEAbhb4bcludlxg/2QBIzeUY7/6dd3+NRqrlItw/c19z6wcUtrG9
ztpz/n3KiPYke9wCBQPa8CUcOG52cpWvGbuiFskJYgHjC+u2W3iLfqDTfaz8toUczPg2HBan2JxK
aH2XwBopYjMTZVlboMunWJ13SoccQru6vm48CP+KrzwyUDGtZEcHBBQIMpW99q/jlYhGxfUK2LJB
MrVgslxl0Atf7bAoyhphrl0TThtqJd+TxlaP0etfk9M5IAM2uU6APkHD6fsIEqAtXiOQtAoohzqt
bGx4+Q3MN4+mzxQbkGUAyJV7Swn0/WrDbDvj/R1YoV0keGOgWmw5ZDADXZazHKpYbNYSuP5YFahr
XZMH+wCIYOD404sIDkLOPz3Lf91Qcbq2qAdzfBctXTQPmQ3/BRTdhAbmFjVvI+gigxJ9zdPqwdDb
NAkJznESxn1xJmN4b06leg5v6FpJFNk1am5GeKUh5OkoDTJU5FxdG711brUz3KymMsRLPt4PiVji
bP97iYXlHZiJ/fsNW1YD0ZU1eTK2pqOMYU2WK5bISZfisJpuxkC7sdPhl8py0FzxQma+apRNbFCq
gGQXM2nyolcSPlsTefJ74Dv1jtUe/8NDgGM9ucKjYzhON2cD0gxumt5PNnoCA2c2AYglnEWKnjSp
JWx90MQ6s6r1TqkupIoXIK8O/c9g6jsOxwxLPcXvzoJ6PsYmVnHOYh531zb/P4vEaSj9UznMC5oz
A9FbswwmKqDbZNwhoUQd1M/F/zCJw7G9Bc/D4OIY+M+R9qOyiPGd64Y7DErNE05swT6rothsT0vl
aUtXt+8gIqWGLfZ85mOG285phvjw4lABsweRadOdXReNN1JK9IxOhsf9q2Vvg+B5d3WChEGmuqYe
G7G2V2rmvcNgiWmt4Y/+EREgQvtrN/mEzWAcJCIQlOOsIAquVHdKSW2Fy+uP9g0xN/h3GBsWtq9r
/zPyRetUatRuTq0fRe3KqY765fjVo4IdX00gOZRIrVYpBumEc2EFq/J/ScF8YbzMa4bUJBPeVfj3
tUrUc14mMCYNemZn54jZgACd+H4wZE9xJEGYvZt/orwmX3utfTfX5DHAa8EcLyEIb4n0RbUtaIiq
Juhn+aPZ1Rji7fmj7yqXQbADfNBYMvQY9+lwWp688Y69EMfDr43H4emc7pPC65Y0TQlUtbwDaffI
7wlyy0pUgzrIY6Fui6e3z+93cFrxZGU0ohL/osrJWKllYVLJheqrQMQhsv+bWRl+uJ8Jvc2Cqu6u
ufRA07B2OdUGP6+oCwQql75WcQ5d4eqZfUxtLCGvcxBUDjwWf9Pc9xwUfurEmsafCTDMba2MV5fk
cD7h/zzOmuV91vcEJRGfIpDHUQFvseAg1G3+CW4vOmfanlerwu9arnygIepL503jHStvJGs/9TM8
nA2QjnbP7FH99f8i9//bx2POyVr7VTz9rtxj9/c8u90tyiPs0qm9KwL+dXYlTOG9aaaUXFfr2F+g
pb/ZOC/dLZJsF3h8KsX/+HYHRok+6oaxvxTbGYNpU9juituSfvvwltamXucP1g3f2xRTxKgUcjlY
vPY2Oyoymdh5MyWoFJ0xYpi4oIpIhOdqewwgSJuEa2fUb+MNcJD2zeVf1zQ1qLsgIuZjOhf4POYL
W/KdDewDSInim0wJLEqhi+nRvJUBRaCCX4JoIPoyg22+ePirMV5T42pi6lZoaYaBiQLBD1DbvQZi
ayduPblDV0hu3txO1Cy73X/cCstp9mu8M0RQ3bJmZnDUwitjFTRU6FiE0Oe2x9NEeYx1HF3hHyI2
1S7IXzDPbMYkvKNTxXvKEF2ItJYDKcBhoWV9IBABaC3Tc1gLsq3HXBgbHhVta4NSS6YIZIzx2m9e
T82CWbDwic8EizrpW+ReF/i9k05MjxySEGmqT1R5UU+oblr46lSctQVAaL3yTsBY8/RZP6pL3m8Q
A8LDKGWc5O3JxLgvtMBGdZgORZZp4NNNmeCfBxuB+AOb+gdlqA1BaOg0cOHh06iWxeDmncYXRWOF
5MYa29LV2n0zx2EbWVDVv20d2k2TrsZAElWc9kkZBsbKFcirH70J8NhOvuKsLay1hqCIm9evefQW
+7fiWWk7jRVBmP1Ip1Oc3c1q/IwLodNJUprbrdgnfiQWrry2adkkDr8rOwSmWYank+nJ6rJeckK6
tvAXz+vBec0R6dFzVn/fshmPplWLLL6IufDLh4Ga1lllS8k8JQ44ZQezKDteuUAiiUK9BQkxdmvH
ugrUsJMU+wnwUMyK280MsHD9ZZhf4YX2G0T4U/H0HPjZ6zdh1PK96YnJmOlgHXO4J84DfiC/yycZ
87dU6ql4pd2kHy6NASSlaNWUei24XYGa8QqsWyq0ESEa5G7slLIXs+AHwcbrjSbFvW0v0zvZCwnB
vnFBDMEepA2xcKnCyJy6Y4OQX83Zg6ICsmikOBbwrwyT856eaghtTqXCSJVEgR9IhFofd7aTEXX8
ZDcakRe4e0A2+34goT1Yb9DFHsvEraOb5nzNOo+8TsS7ir/ed7qU5f1PAB6hqMChn3WvTXQvl/Yc
li1KEMhsxfiZ3HlYPpOpjbAyeZfCi2L9tF4wI6St8Ijx4O/vOAvBAZVwD5wl9lYh1tUSGnNcct7O
0HwYzr/J5D2TrUpd/otevsljLytIGkwyvEWkBy3YQ7Ui3u7OGyf/APbAv+Fh8iMCX2ZN/I90DcTj
77AHl4KkryIlg4nRC2NNAUoxiLDYkriqTG8n2mUwY/q2DgT/UceedMw2nQK7tVIEgJ/I4KGUlwXr
MXsX5x0qUh27UCvR8W516d8QRptbvlMIPN0LMPlVcr0UGq4ucyfHS9Cbd8+miFeuwBBwIitUAWGG
mjrXugQG1CN86MrCxiQvPTP7HWTEi5Qc5WbE9UdTv0fXgMsYQyT2RjQt9U22pJrNKPj2op/GQIKj
LewHErJubqNQc2ZiMLRwlvvL2gqGVaM98PfTdIM8m3Tu/Zb+GDxElK/sjfVD2XJj7VNX9Eewkln5
JJ4iXom4vb+Zk4VuVbOXYN0ixmC3t8pOvPch0DVAW51DaHevhuxlX+qCCmepvrGih/YWpNA1nenP
qYq7HN25aMc=
`protect end_protected
