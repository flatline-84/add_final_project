-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
sO5zbVnZ7zuj6p17z46JqjLmHSAV6FRJ448DFL3aHYugZDScePbDF5a0hQggVXB6WKFRd5XVAX0n
9BE39hHZPpm6DO4eD9e/3wuEAnTC4LwHHq6D7A81ky0sojmqXP5aHjN5P/w4ktxPPT8gLLuxSj0+
DsoVNRVN5PFR3ICvwOXHwBNGdiEu3hqGZr+uY9rRNz1lp1chli2M0fzj7jC+H1Ru1sIdMmkrW4nW
fmPjZCXJXT/y5ZCl2CVYl4b5AhcnTJGAvhfpuYbXpPDOk0n5nB4XER4RM83F+9zkQigifQ8x+qf4
bIxt7yn1D/tM+8iRSBjjE6ncS9PCwiEmWKtEbQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28736)
`protect data_block
AC6z1w3y6yZEqM/URUcC+zutVMsj/xAJfLV1ZOHLoAVHRaUJkhBOB1SIOFGrhGaerGfAk04EzC0/
iGNsDm+Pgui4an6WewoWngvXqpxHGuToGY24mMIfX5Nbj49sPyhvlXrRoFhfY8VAdl4BcDlGmFu6
U/3+2ZINLBi/Oqwdmr3ma5BNvs8ZXc3qHKR+rFx+5DGSOqWQZ2TPOfgMrsg3ljH8Yt7iado6/Wed
iM65zGFk03kQ/QI04LCKbhyb0NHitYZER04QrYSVTNsoCME7r4vkR+Nl8x3BDEfWbBf9DQDClFdR
VgOVRwpdAe7seX3FIKr4Hq9q5sDSFD/ivt6A+gGFupDR5GhvjLz0WdETIO6rTPmaUnXpebNcx8zF
1o1R8QKrfvnubDUkEPoq1Yg0CeavAGt8r550rNfFSA63eQAaUgse09p4bfS/L/1hdesF/2ZbCZDS
kJZzBZnV9aXq53Ws0G7CRyKOfFyD3lSsO8C3+DiYzMqdHDqTBsXsqe1reAxMxdtha1aU26T/iJeu
iMvsPBf5PrhNfrsPrSppf/7Stm0UWayd1ZxniWlgZNE09ZfHKw/yRlHjeyt1MKE+V02TTIoLdem3
QR5yK/J9CMTFOyVBuG0oSussdEcc315PRuv4p/QxKPComtFEK3T/r51d5jR0TG1USK7TxbtINdpq
eyR0Y3MANQ9OCG84/4RvBzL+n3Js6sfVZKySVYbvClFN5kcfe28DVSpySkFj2ESVGvFNSLzSIfQm
IWUBVvR3+pnYO6C6jgyGLZRjTOOLaRI0Tw+zNajftPoQrKWPcqAQ6Xiu47BL8gHH8AYne1+tmc7C
4fX/TR/BW6EcvbrkoYT5Erz5q6AOYpxgxShiS/TGocO4f7n9TFyBAw9UMBiq3XWlOn4ASFMdINvn
d6HMwS/mgM7Z11ED5wlHQPi9bpwpYeI5zmoO9/li+AZfB9R3vxTHLaFO1hNt1ybxm11cHJx/InEA
+/Ht4iFZoM9BUa8MtANkovrgUxA5q7IKxZIdzwWI7DwbFEmtCX9YC3FkbbAoOc0uPbWUmO35nPzv
YGhPp2baWO4IVDGM7FZqMswYy7rMEAuqlOKjqkfd7oJ5GnxASoExPzOHIGgTpvZ4ydoooTb80kXJ
Ci5q+C/ZypEf8aY4kAgFlYxx5Rv6vBYgkkf6Eh5jMtPhaH1OmYJA7PR7UmzH0eLG4rvpXEeWWyO6
Fa36F5HL8a4SGcHdP+OvUARceRuERdY/C99o1kyFpw5Oeeu7IXLcRCk2y8ICe+wg3hpei2sOc1O/
yK0M2Q2tTcR/5dwLwHNrFGzQwPekvTxVlxCzuYr138mj9EfyU3Pd+XjJTnxishUym7KeuM2zNQu4
ZOw78WVc4OkWyzNbfmdiQ6pSfocfUxW6HFtI9vlN2yvyjeR+ZldfbL4QrjSMIbiLetfiymKAVPG6
elvlij/clkpj1ZXo2k0i2BG3ctrvL9hBWj4E09NOofjv9AcDqqVdBdnNXHO97zmUgL9h+uXmMWdA
XLPteMloi2JgqrVHxbBgOV842kHHLkaI1k0ZkisNiQpNdbjhYJevnmUKk+ePK9FdKT2epA5pI8WM
xisv0v576jluhTp6bdyX/BUfow6emtAcUGCSVbv8RmIR+IynWaH7TAL92i/GTXrUhy6Xc8hAcugX
1bQHEHhgN7W3MWyDUCLnXnf00kSCa7ZJIp3LLagWw2AuvkRHipXk2dkj/9bVHoD77HbVd0/IoCpH
sLle25WhbG0NphgRnQZQAJU+mZxo1/7st8BxazGrw5lWYpoelgNdRIkESa4xxSRcAT70Kk+/AYB/
sNhS6njivsHt3K6Rwtcdyb93RDogcx3o0ntkVFdx33owUNkeedkDeEZpTHeeA5m6q8kBPfBK9Jes
xMh9dTDWihP//2x/do7LzvMOeo6rROKUXl2x8929ke5Ocv6PUoH/WGv8KBIv/idUMJp6XeNCiF25
7tGMfW06Zw5eQ3iHyTdFbk6JbhkoiPHX4eaF1OGvxfn1QNC8kKQ4dx61dWydUiHvvLXnPhfZXEg4
YOtHv9qQHoiMCWAwdKnckAmS1eBQfcJZ/uJax0UEElrdcncTFozeGkj5ea/4NJ6yKTLGGwwaFX3Q
sZyAc96kZpAJwmcJwqlwiJC+DKofosInt++XoAUsGN59MIijJdyhsk8J69ejCJd5WhMNXweSXMc9
DQOx8N/9u5mAyfVQIGbqO40PqjiceD0sOpCALeNG5sW6FC/6E2SzmV+fKFdXbeGRKhGoPcJ+osUF
PZcVBbVmIJzErqfmFQ6cX01NV3u9yQt1KO4QgUrRaUbteLtR8b+t+Gq1P9n8411ITMQ9ujG8/8r8
wsmV1rpssBVeS6yW82bgIPXiKyYcmwWXwBi5sZsg4d7pGfXgYX6qtY3cWdAO5piXjdahCieb9wdQ
MrFRSDv0wJ76SPSH60Cr75Rx7gSXwLO9ZAZTTfi89WB/oFpS+JK7V3CzS9/ybDNlK6mT2Oa/nutG
snxJFiCNkLiIgyOQP4BV5mQFAZHN5ds+SGLXj2UYXKB41Q17Aesgvx5RPOCoqssn3KhzapJSS1/X
9del1JUX1GzXsw2GHLbLu30rTUuUwvN5TlSjik7u1McjCZVuOBeAz3nJPLrDaMr91go8xVJlm5WM
q7+KwL4Pcb22X5R0F8HwoWOXj8baIbcwooSPtBoPKEEu/k3Py2C4lPiZmanAMBUagCn8dkZx8wz0
TqL5bpd55RoOp7ZZTcTqAxFiqUWEja5CPlcUVIgVT3Q329odBtj047rWAjClW7xC18e9aLbgDt6Z
3rAkUHxHhYY5PTeoYu62Id1/FhR/XazDt28JzODTZ5oBPImNG788BcKrcDAjXhnwF+UdEzb0eAY9
8o+C/m2Uf/1OcxOBZn6sE7irjZ7q/KoVPxEC7p1DrdpAjERADyt7SzyGyzA24ZqIzWVUecTwdLAq
CdUM+lOgf+KgY6cdAosS8Z7ii7iBoP3cnTLMzwE9ls1xmwCQW+v9mk3k2NHADLKcLDb7p/2h/2nP
BK4avrnoVb6x6eicv/WOSnebhDl3vp1wcgVCKjxqVto/XtHJ3e7nbk+xNZ1mlF+WUzvlrC5Qn0v2
mfucLBP3Buxn0m+eQHPQDLlKnl14J5ZhNO51PbrcvpVyttn6naQR99rZNLCBowv2oEqi2f+saUoG
oazhEoEj98t8Z7iInggNa4tCpIXDIEZA1zLiQlwG408apWz9QJF8b/ZIEy+lG76j/MTEXUV9mQQC
iyFmFdK+YWr+JNKvyPxd8GGYEnQAZfUEbrUQUn5f1c1vSUxjVFNvVvaci/jQaQmm6/hIxeO6sJTR
OPHyvz3BKab4AYyEvsSybZk2HVqzLSXWzEr6dGaEJj+TRjdiiCYqR1Yw0uqToE920nf0Wun/kMkI
AiSuh2An149qDV5iFbdnBsOCXXETtD/7WMzm32XiWJ/LvS8MELTqUpdCgNg/t4oQYRlpDRJ0xHi9
TmwFA8elZQOg81vLvHfCgE7xsVQoIssDbI6MXjdPydMeWvmaH2G9NK3CHSe8Y232R2hAnEiQkkS7
qcfu0fRctb5uGJd5aKoGJcBwyIu0Wh/pkt7YNR/3IsMpu5f28dtc20TfP8npfnkk1La/I7beGCXC
lV5RlwGFPsOpCj6/8pscsKztS86jSDLDMKngOE0Ev9h66sdchxirqJJaG3wu89eu139e5p1GDvGZ
JC4F81NnG8EpL+D24DDqAsIyRYrRRYlPiFBjozr6d6lgIBzyyfpfIfTrMPjNrQDRKaRxNlTEdD8m
9TDyyAWRTmT/mosBfM8tIgVTYzk6FbPj8UQuetDw3oHzZR9eZt33AqkfNuVVDpVcVGqoe15ABqU1
P31uc27Coh3YinXbrr4B4lg7Lx4WN2WX9Iz30OWJQtzTmdqn1tgIP3B17ENg+emWpQj55Zj0L5h8
yA8nwP8602FUkn+dTeHPyGkR4+AUCjy1qrn3KjKATooSrLeA7RuSatreXvX0PzBbfIsm0Xz7lPD9
UY6ycML+C81mVRFGTTYDUdcoSuLO1P8ZGQ8vUkBu6rvJ0sbERcnjinG32UBa9yfoGUtSWAOQ1UmV
3J3BZn8lQrvOhdtoes5LE3oXzicI567ohU1dB8PmLwhWbYPzXN4oXrSwpDZw+H9+W+avOTvt3rgz
bRRvDe3rN2TFhCOJ6ojagvg30dMxt9rkcDAqbAwDi2EoFr9ioYJ9Pm1ymI6OJYuU7oDwVeDQOAAr
ZOUTDIef4CZ+crbA53m6uOOzFD3JfvWFcWIHe5Vak3RZ/isXo3sePQsBCUJk6cuTyeHNthjivBuH
6LJfCkrSiIZxFE277KWFrHlwE/ZeUrSfnQ/vBvXgab+e1JvOQmr3Kra3OuIDAJUOTcqy1jGbHCZJ
GCWMdfWJM2zZ/nhYINvjyIstkrBrmq70yhUwReeCovz2438Y/ZZaaAbeJCQvsLW3wk0NAPvoBHvp
1yjQw2v8KscAVhY4H6peHpyJNZQskdelLKv4qtSWpnYHNL/JM+KrFxXIQxj4GRERzeTvOpA9xZQ8
C1YiaHXpqxNS3YBZxH+fwgSb9JVRFTIaY6GH8P6qn2Jb+GR94upVixhT86ih+DG5A81XvMcM+nJv
rsjEZW1QySDxx3ebF95wKXZ60rKyqpAA/mAq5fVyhRyX1LMTv4LL8j3EoYyLSJDe/XqpUQCVwUK+
MmvXZwDN2RDI1hEb+4dnncKHsPXYuYb7COzHDTSv+8jIvkfLurY9mmoLqxB0bG1M4++cPXk5K/gz
b99pWo9pDzNhBaOmFYNOpUJWs6+pYXp5wccHP73phvxAByaNawlzLynfP/lKZX5W9wteSS8cr0+K
NmfgvVJZh/2u+aKQGgdPtIBe+4xmGmHCcazaJveBMGN6KSdZ47ANhjCNz+NZ7yFRbIqvCAf722fO
A/fXUYHQwxvrrQVfnwoS2iMtGAr80tLeIHCKp/vq9fYNM6Suq/crzcMBIkOwtGINakZDOgXt6E5k
MxinirTOJGGxgDixG+XnG70fbJ8FqiWH4t4Z0qu7JZ87vK0DQ18jN+m2cwK29G8FlDWLEYctwRE9
SvHgKxLT8JdqpYsuvI8Om1CjC+gn0BtNbgkiHHPOxqQd3ElB92GQidEhSBeDhihHWUnzrVwnotKq
ucZUtqjtKrP/xGSDmZ1uA8JwMVppLe4CzAVYcbbm6EOTjt60eXu9unOrKZSrPEhOA5tn4z47jfoT
QzsLUTU3IreeKsvyVR0aGchY4A3xHOdM3q5sFai0tMZOSkF04Tiqe0rPkprZOe0HaodwEJluZYi7
IxsBDkU4/29u4ioGE1a+m8/JZ3+SJ2giOKocaHbRFvoucGPswddR/Q57n2eLVcw8GjqACBkkkPbF
8KYfoR0qpAsehmDuVjuofHEU253Cezh6G0A66MYI19Cy2WkBWmlqmhe45b9fXNhcJM4ijgY0v9gG
0FAn8B5WIhrNYDfgs1aCwnXjOwUXOe8zxKiD1aBtLv37qUkirOkiOyp5wqEJQSaM2cGYOfAQZAMa
1bEG02ddpN7jILkdQAtlKbIJEq9wDLuzaCMFhj7DDq4EZMd50GtDhnJzJy+N2FL/4wW1MgrAt6ah
C/8+OL1qQ6XP8XmpfLe33u4mC6poim8h5PxJuxh6vOdcy01mZ+lUvZKlMlvY/duYWHbs3v9hnjOd
IUIvK8Lq2Ut0TO2SdEzJFc4Mux/cXA+AjH3zeVf31XiLikjDE7+Pu/WU55/FcEeNN163XX9J0hCX
vr4RqPTwgh8pw5zlqRuq3Ihy1jVCeYMXPwbKdnXK25SRxnbqO2hq3JiIMF96iEuuOMX/SOEbWsF+
uqGkisHC/HfP6jRYAM6Pou+09PuMqpAIb2WVO7Alb7LWK7LvOxjO6dP84aPXjI38ucguZ6kA4g5i
0lmNu46EGooksDhvqu4gMRhrXQ16WJtislbBBbl9mj4Jp8iLavraENbAhYTPzjhgf+KzVJdr1ccB
LinOZ/y2OdCXdIlmjVQBABUBc9Qw/m3/JRPqxUlATsrTSNo0DuiiEEKGfeCQl0t54+sBQCIEH9x0
Ckp59Nkjuh/O3Dy8fv//0PyvUWN/f7HnWqMpCNjXzikjCbVqBFNkhPYsRU16x2LQGa7Hb/OCJ9yd
Tk+nI9oG8s7ES9kdVrl8NAn0OnONAAo5mnW41WQGBI0FTTmLDkDvkvn+Mj28hZWsuX4BulU8ygyU
Lxxj+aTrT8cRmreNexqP47Qe6U8YLO+iTEU+nvpsZ698N9OPlGSVNvDjR4JzPdiIzjV9Q3B1gRpY
lP2L0L57k3hNGijV2SobTeFvkk3M4xVCsLh/LYLtMCpS2Ukt/BMnJS9kL1pPfVfSLW0AssjGZSe5
E154hPVQL7bEgTdFr4hpXXnfKm1aR1zRKRA5KtsC10UVTJLGuwbwzm+zFsE34yGrhPZFs1bCULhG
70zk1UOJIzsQPx3pu05piQvodKe+udLvOfr2Tt76uOugNx9sBE0FfOebPMI8DxXOwam1CmJdKNqJ
frDk7FFXhrRcLasp8Q2/TBhMMQNerZLmHmrw61s/r834zm05pORfYQQ+lW5dOekfen60wvl9Ivyn
4pDKDI74u2Sob87UFKKELXOEePsDrFXX1ZWZ8BUwf4dAf66yis6L8y5Cnl+vn0Z5HX7iP/VunZ+a
Hfv8ZLrQBxtTYWniixzclenbPe+FAv1CDpk4Z1gqfXC8bXJSGGEB2QfZNGbS2XMbs4l/IDe17vhl
1RDddO+18VGkvCTBW4RrknRvpc2PHMzqyJL4cNbeKVzpE+4zLHUx2BAooZkHG1z3H4H3AzCxAtgn
cmNsAE4Ay76KPCx6TKSUGOnJ3ZPnowp40CTFW0nUaMznmMlxtcwlstItjiV6z+U7OjC8/POjvopz
G8HuI9dH6ye4+yiacoImSI2E03Nkl/dd0xiKh/MCmI9DUF6Mk6hwKfU0LGptnxdFSdOxlkKI8upv
LI6kDc0FHdoLWoBz/QfDj2BZDAi1lpHGO3n+KplNxAe7bFDd6FYRy3vOuNQst6aBW1E8TsyTf59R
IqzrVeyRomIUYcCJkPPcqL7uQc4wKtupP97EZTUjIPwhyqB0DTHaaTeQ1JQGAYT2wiC98mnE8lFn
hPA81bAqPBBnrs/viAX4YW4if9qcXLGN09gLj9I3fQz/Ae8kxiY6Dc6+NCU33ISg5/daa3UjXnE7
Z2Pg1M3jgypYrMAHOM3mX4eiso/aKGZsU0hCzVD25G0Ukr4rvi988L0dHo3etbnJeT208OwfLcvc
btN2il6JME1pCJCJbR0iAekLsbf1LPu9EFkjAko8gw0LytgSYqvw4FQ9VKqkbvYssuVUHNMkyooc
z4ndiqoaRCNqtjsz/Aq5SCfHJ2HRFpHOKYgtVHhFrzjxZxODhNjjqu5AZmQRXVjdumC9T8xX0AxL
6YZHaGTSzvdKoJ5y6QhwilCKki74i6y7ktRle2u8ClWewk5EzzWqDCDz8q9mhIegp64SPCYhDgdY
S6qeIs+J+v1QWUi3fHwx7n3ED6tx8WTPmsUSK3GfjrtLyr3ZUUM/tFDUl6OtRYZI4uhgE+UT9T1u
4cTIuXxkPvLPPzPNCyPfN4FvBHhAvnfolk+mL8mPvDc3Dn9vCVdQifOCDQgcw0zFhiAsjw/I2qoH
QfWMtbZYALFSG0KHpfP6It9W0Z1oM7qopHrowWWWl3y8d2k0WlwEX+FWVm+gfgWtiX1EvlWkev68
OY0yShgvU8iLM5NSbwpRFDNXWkcQUetmeqH9axdPF9GdoIcqKU/rGY+dINRPw3EErnyuuG0HNwOl
clP73PKz1W5WS69BLMuK9sSt//MymZTJCvfaICLzXcIZJXDM0HsmHG9kkwZsUBrzFyGdrEejLNIP
F7jZYKiQ5LuDnjZtasdgcVSSLnbOQHjNpxj9yKTIUGxoZ2XEJBpGiLDl0NouavIi+E3M5OsMhlnx
7ZmjuYDNsdEsAU1L+SFt0eSwx75m7mDsrVCeE3kR1Rf3Zcq2mszcWK9DuUspMEDE9Io8OEiC1G3j
c0+dBglRvRxHpxaJ2WsYl54KY5KC8ZE/xawRi619jqDqO3v5DboDVgfHVQR6riLeNk542zo+joOZ
Hun1yOZ/KN3GwRFXOKvcihcIzoA2flthHE0x4p5fdCNajzFbaKy8B8Odr42FP9Rj5nJfbBAydxpv
sEG4MFL2a3lL/bd7GQHI5lfCxlbYXb3VFqG+MJDkdQZdmhVK76AeyMdz1w+PPBMRzUtSAsgJRstD
ntzNkUf1nvWqjq8LYU6nLoF+/5ZmfoKV8X65PGSJbQQJW9BvjsfJYsi5EUTxmyZcLlczPcY5k18y
rXzu6WdWa/+ldkfGZIkFA5P6dfApbAKUkQlEVffVfrgLQzEvJ68BAj0Wj4pwWjbToa2QijKs61lR
TJZviiWBCDg94bPDf/qlq56pr9oGKPq9XeOp+A0u5mF878eVRFnIOwF6RV9bTtX9cyqIsX+oF4rh
dnDfEtdBARkocLOZt8DdAawpXgYB3Y2CkErvtavpIb5UslOlx+ZNAtp+zzyz/W1PFAjsNOqPlnb8
Kl9vEtzJQrmDIhV9iVqF5YylGbqp8uzhRblCIcSvvwWKr395fZtGaKY8xnVBrrK6G4uCohkZQqPF
wt4fElwfax0I4iOknrwhO3X7m/08h+0MamIva3BshK8uDAccxO7gPAAeAt37vNDu+EQljinBN53E
7FoeIA/q7MbaPfyRhXoWzwyXk/1gD0yFPAszD8C7QXP9W0YZh3ApS1qG7Gf3PvlXFNM9V6dUu6+N
kOIdr77KpDLxjMIQCD4NtWRIwdHOjaNlYPggICmiIrD4xFOL70i6hjXwdZa1hZgobCSbs4Foxq0X
FRrCxY+ctLWcP3rR63qLx1y8Lf3fT19KqfNDKmjd9oSiaMiOKqONPLfChpEkAGd9Apv6J4QaMXV0
TAjB5f2zQJjI5klQ4vdI/iF6JLWsuO2k3L/PaQPWsAoGfKwO24jRX+1EySSAPE6pCOGLLsZB2kTP
WTQWH0ovxrR/5eq4IIxAV8nmg6lTJWnqFetfOOvtuKf06j3HM/VaC0oIp0MzfOY2TRFqGFcKmU0m
EjpDV9ZcU/yQ99Bnae76CRWBP9VM87pGrRk0ZHcEzwpoEnPh9wkg3zYInhMudfkg1D+w6jFxpj/+
o1bHVjPRtxIAXmsNUBgbWByVritjsvhJ8ffnQgjiDLVP1qCQfF60TY4cbtVZLWmYn2lmp2vEN8Od
sm4hZhrnAf25JsgTB6+1my5Jc9Uy+rimUrV98Zql93zvkZDkwOS6hbtAAO0HD3STANiagaY2VWjG
/eSB6q00xe+zi9gOU3WFfGyqs5PlYv/1IMWXYqSCYr7IAkYmqCrnSHPer4pLcvjPagQ06upSLshi
OcmnvrURe5bXQ4VBvHFAsLrnZI2hhJBebg+5jroorR8g4Y1V9veb4sbGsELO0R0odEYFOBPKWGkZ
tMDrQqqQkOHKnzxXSMyHZFI8blpwp0wUWFrXf4kiPiPePLcieSK0hgDBrxeGgAd47bsUYBqDibsg
mg1ZLcqnTZNNYdS/DghVh+0iOHdz9sJcC58GAyw8KVGaDMsWi/sUiC+4HHQklvi2Oa2jwc6IYQgF
f4MXvLEbQ9xAdgw7FmG02/KLZdMxAdBqYKDt2nkUnPu7DYeuI6DpGHLwc/4RZtA61Iv/3PwS/jUv
5JA1kCZ0zBG2j9gyTC8MWAoobxOfLX8aJhFf2gJuK4BTV9y01fvwtCytLYDCkHWZh/XIjYFvVd0+
kOEiEXP2ZQEifPmDZYMs8J+Ek1StJyL+QE40JUlNjukRfbobPFmjsG+ge5pkPlU2upZLPxkZS/q/
2KGoDv8RvIgrnifbMmXCaAfOR1f2KqB68OFHmF3ro4EJBmYzrlPnsh9amlJaArT58mBK9irWsgGg
knMtk5PQ5Z5JUJzrxu9ja4FmVZobYO9RRn9ZeBR1Qh1Eg2eRmYYuU6NVuJg+i2PzZ4wDwkHOl3Tt
Lo+D0dQaWi9Ssq+iAMxtNQNKEcYTeNlU65HTnCaRODPUWoS6v+BMp5ihRC9s/VHcch35ajehw2on
Ugr9bgVJkP63PZPKptYfGk3w2VaPvrL+uAxncvtumKvIZYGs57DitzzwwcrKq8ukQyMHhpSv6eYg
H21HvJact07jCJP/vY3zqJSfm43aW0l+q4Czrutwe48B+hkYjJrhK69ww6WndcuObpskNcoPr9j+
DNhjgULIU9At7V1pN6qa/r4iSRBpr0Q9st4JbdOBJWLQpr2KzhthNI2zjUXBIUBsIX4ECueVSyDP
na0BYLC6ptXo8SFsmiCXnj+of+5MOvOq40WDI3cp4Pqari5QodWj/8ETv11f1Bij3Jrmo3Rp+CqP
MYkfv70V93hGf9Inw7tCELYjYEcfua0BRyXMktILgY3qN5WGtzqLuRgn8nAWgX5whKsdUzLpvZvx
0QmIXnEykn8BrjocYSTymtbeKt82fF1bwBphKO1Uea3ftNHOPhCMMEAXZt5sbzsC+fVZMDqsajMG
OOsWHLVPGi5oASE5bqtTwtB/xhUQLJZtO/IkpxCBORqLElH4pODvS2cMYeFdWCl52gkAawRJsh9z
u1XWxuyxfhhCWSKcKWrA9tbTuQotqBXBVoXFpPdmbB9SKG6e5a7LSlwQRu3dDzdD0omOfo907Qiy
OV9KtEoGBMg9zmRtoUEWkn2d6pRA2iSyU15nIvuEqGSRzgrvXaYuzpXOgTh6V0cKmMrW+ETRXTFD
q1IU558nCldVY+baOLHBnBtgT6rqfolwlXXYX7qhX1au5QyMU8Su3wy9IOy6KCEpK3v3ddwsGkO8
2wvFQquqJfabNC45lNSlFLzhnpmcnokE+0Ap1wjG8dnwHyTuYm7tJSTbsWonpYfXqGp4iR9vyju4
EQWECAmkcGJg8+yVn3NgmGX2NmGVTh9H0ZkUdo2Mhq+4VeQkUvFJE8xqHwoa5PKCjHzhNuPMuA8t
1IrJSBUZBzbW+IfOJ9ZSJIbuJODTBQ0bqCXaeikpcLAlvfQBYc03K8w39t0kEVVCgr/xfRKVcLxq
1psdmJSAFS0qe/vP8NchoMmF/O0CJFXB0ewH74U5ArHrMa5v5Saa0FnPCMC7gpA1RBxuwmqFjtEc
SMFXgzVR3pJdPx2PnUfufj7DJlVfNWVEs0i5Ns84aulUkTP3zJ6bkX9TWuUE5rL4geo5D8VdiNHS
b2l38dvf2zHC64itOHnE2pN2Ttdoxaf5y+jBiVNboA3NUyE0ZMJ+w5hdWDQXhsV5GtGrVczJFC+d
sUqjnL/9Qc2T8jeMeF67xDm4PxzmM1Pe3lsCuLGotV4GYzkf3KR84+vuCg5Rbma2MX4aU26wMbw9
Ved/+HozkZ/Zt1mLz34I9VizJOnYx0s4L/AjGp2i4qqOfhTcRRQbvnbxccFIKArz1ijqGkoe5+7C
LQom3sfRAKo9PVHFlE6OT1EJ9A257OQ8zaygeGqeYUxaRQuC38t37oD9gp2cSC7zsG64XJAmwLDg
MgRJkKKR8w1AbDsLFFc2o6aQ3l1jpJjGu5XLUWj6t5wunQQ15o3WU21pHFSeaJzgHzo4/JyIX0Ww
FIVV6hSI7rPhQeTIrvzTt/jtygaGM1yrugJvWHbzszTAZjlHEidCPFrILeXzU+lJ4ifiPrn2ybty
2++x2WM55GJJvR2oeGHXst1CxcKJpGxOQCEx4as71FZliXQZawbV6xTTcQN45/ngWYZpa6qpDGDh
NFFW1adpYjf0fhIOZFQVx/T43/vp0HAUs1t9mmNTQ8POb2aIRFW/XhLaH81/gAAU6HkoIdUkNVky
gKK8MX1D7tjI/VljF5/L6x/6oEpDvzJdzUheXkLb/WOKgzrix/QK6RIgyT7EKlSlC8UBrD5oeJ8S
6NcXqp4Ei4Yl0Vu7QLmi7UBjXNP5JT+Hf10WAXhmPH/smVeBqfQhUUwPoCEB+tsfMadmQVtlcs+1
WhH8dy85kv6/rTvM7b8bncT0ZU1DEI/YDVgImAmUba6AqRm5UJUp8Uze9O/HOYqfQ5Ow8CxejV3v
xkejsxSlucLPcMi8kIYQVggEb3oyKUL0CCdbhkNJ7lQXnSx/S/y7wMAMSMFoUrXMRT6kSZEHEKCb
cAwdxl3jmqYRP9hGzsEfcUOjPKq8wC+xwx4QEpzh7hyeAHZnMrq+zaEXE8vqlNRaVS9YNIqRdaKd
xfL3byhlLHf25p7lW98A04kZu+Yj9JldgL1bFLE6DtLPCuxTIoO1FkUfBIIcDtL0wLui4pdBGiuA
245lbWHr1TqqSlpDi/V4WsHqN1JmlG7mueNRiY29acrJ37e8+JknFmv9zZCEBtLjBDa1/q3iBsto
wuWUzcfh6supfOY9NrK245roJx12QtQyQUvEhL3oisgehUWPNIwtlkxTPxRqorC9yO4Tz9KEW0iq
ru0H6vRWLIIthjbQkYqAnm08YrKJ0q6VsP8RbSESmkTR5iEMCkOsdMUWI3QPPm/0ufl3pLtWe1LN
8zQrawKvDUHr61qGeqNZZTE1U0tZ5R0gKE7knMkynXkyZm6ngOmV2h8iEj9diGQp8lubROR0OaOV
bn2p8tXQ1qoYtBvocPwmUo4Eh9yiaxmPTVmPDV9k4tirLEifcKg1/mp83HAQWPoqJW/yYr8YaGjr
x4kjNy9Ipqjr/hbL9fd3xa8OEZsMSIJsdxuwyFtDBbZA9pVRbIybqIvTNU5BM/Ts1biTNKQRG6ZB
zI86uzTdJm8FR753WKi0yGYKl+I8f+ZJ/0L2UdT/ien65iWoQjzI5KJB6OQaul42re7lMTSjvji7
ScNmrbgEasmUHUN4Pv5nVEqmNDFttW+HxExun/4ta6Sb0parV/r5frArSPjkJQbpJDiHeAuRsMte
B7MyuNjk+nECP/TnkC6XviyZO8QSh8MAMlGTqXCTujODdM0U6WtlgpKQEumjFSyU0vouivOMqH8b
LgbWinh5un+VWIlpuNgjnNwSV0mJHu2aHNRmC15Fn6/knSVTeNadpz7WclwPi7B+Y4gvHbQGFaDj
SuBLLSnZhO6x5175I0BEKd63WcjaAgSb58noWoPXSDLO1dRrqNe6WL3hqqs4iJ0wziMPduxLRr37
fxn0r9Z2CbIQlQNk//7HrDv3m9a1W4iazbCLCGpBcrran56MQTEneLc1vWD4MJz/lZD2Lu6Pgi2/
776D6sqpr/p9p8UJ5qFs4y+d5LbevR5cb3N7EWMPCZe+OQCZ1zfewH68b+eOWCwEn86VSp8+pVsQ
o+mvi4cZPPJ8EzOJcz4vYO4w+1q2uIKs6pTjDH548jAzv9FupWn4KHos5EviKQkVrpHXQweeigjy
PDryUOZ2PhnjZjwNi2r5/vqo+WKeGB7TRWr+ETHYyeQHojQGaiXQN6L+BTiZI6OXeFvh4k/ENR42
fz9E8yxdb9fxfx/lrrdV73OmSm256ZjQXCPgMkFZW9CqphsfbBoy12bQeqUr0pgpwtYq6w7pu2dt
bFsLtNaDwjgsp/duTX8IPM6GOVqpQVowaA4bLeNur2dng+/Q77WRWKvNAT3L0Mj1p+Hv5nU92IzH
menpJVUMuv5U6zt9WIwrGkUy4sk+DtLvJc1d4SiLz0mUT5FnZpoVGpNyabReesAqM4sQPDRaZR3U
9sgEAQD4VQcc19s3k7fq+CyE9c7fBM2UCX7dXUmCGhGSLHR3PTrXMqwqq7L5S5p1/uC708vLsmJZ
3n9KDH4WFmlJfgD2TLuSd6Vs65zxYZyLZ2XvAa0VYPX3yJhfAYLXSyYvJns1kavW5EPE8JvTJ5gK
QX0GYzlkC/cZO7ufB4feZgC5AKo45vGFX/k61CrEi1wCwrGud6ekNr4lJtEHTEGXjJRFr32n6pGO
OpDBy3T2Tqx+0sCBtS9gnfdk4MSPfKBpaWeXHZAJoPY8PDv/3H6F2kOrwrt4IoGhkxQHm+tUnvfV
oG80Nl34RQdbf3Kam/R5vXUOsXEH5zLieMa25VeYBKLRVsmR/gHLDs1UZzeD/ZG2uoQYfEWHhrjB
0ThVHgGKqx5DRMxWmcGlSLW+3Z2lEzMtErVb6kgZNCi7OO5YzPk4x/Ypm/5uOt042yINJSDEF6nh
K5LEp93TRIlCKFTzAlAy3KXbACIvh4qGFxFtS4oyPBCvMWgCkuUTlB24MtuiLuDag7qhUMVa19T1
oLE1IMbDrQ1U67S6YYnZWho7jepWtQzXB1dODiMNyZ9PwlgIAvCn0VM9idreYlRt+a/zSi+90jX7
PVxOuwO+VMqq6rRRBaXxSBCbjkSJq+yC0kIX3Umh4wBmTavLZaToUBdAPGsrFi7mz4CO6n9OxL3S
eqBrN9XUGBeyIfdZWhniGDxz9O4rELJQuH38agTDe0Epk28j6EwDg+NZhl2cJRQzCmqIiFGZ5yH8
coEfrJBt66EOghbmRTbyVQaVmRDDK7ZwrPto/F9EX7VKcAueanlMnvuge6dhINcA8DTt23ZZqlIq
nWbChq0yGewn0LMjTG5YYicEQRLeqHLHQ9T2gZ9MTTNX3RMkKTlddU+bL5F0BZxRChxiBVrT+YRD
pRb5tN1zE7S86+ykY2a6C+UTiJXXnrQ+CZ7owe3ylNQ4flBVCJiifNHZvEznkgTEwm77sE0rfOAt
90dtV6ZDjt6kJrlxABmUXwp3iRBtc3PNZraMokHGLn4vi5RArq0Jv8Qff8+ritZZtoxUhV02eCVm
Mi0uUltcsCUBADlffNe04uebCoMIKEvZwDakn7Mpyt6CdrYQaiAPPtILlN88wd7SQyMVwoC8Xojv
J37Ymx2ujpw2FhzQlo27kAagCBDaPZpLXzXGMPseQG8VlhHPncAraiAwUR7IPaPXbT3T0OI80twy
gGyx/3MF/aUGMKG9RrzY+kmENNCbaKszuaxNcL/42q2PvQnIORyc9s12+CN3+EU9M/NriRmLWP1K
ollrdJh1mlATHB3YIVWskvqSgvddMhhjJtmq8xX9fGEDEewqFT+Nnt4xDy/GlbvRl8xTGVq6gWP/
xCIWhAsvd6FNV6YKJ31ihn/sPv9twGZsJ3WBYi9vI69wIUI4EP0P7jhBfH/GpoUw+4AnuRbaw+Sn
e7SOKEfhpJBu+tPSj5hXoctpkRxwh5nQhYJ8DI1BEw+A0o6zLYTZbsThrV8T5/dd+UBjjcHKFLYC
7lnOrWP5rKBlUjdTqctiURRTcVSWDPN1e5UXe3AibQ+JvK3B2QlXgrKhz++4EKR+mkdosrKWw2Uk
uyrVcfX008tlb1uY6+idB+FXCqF1YdwLO9eLXtXLsrP80617N5ZiZFIOA5QveaYPicIJg5cmSRxo
Iu7ypoRZpw+thPdNFk7iJG8wF2hUsqgrBIHOyO50fm+8+M4AzMd88o0khCVtDmAdeujSfLkadu7b
yXSd6snOok7/k+VZPiSglubJBXBB0voE3uieCVKO2gn2Av5FSsQTjoVl5oIppRNNBEbQ0EpupwNE
KzoltkV2bQ6M+4ejh4sY64g7XawZsEBqPJ5rKR1mx15HX/vsCrbMSRWrlVhdm1qT9eQOSoKdcKE8
skzWXRqBL7wr7Xw2m05rCdUYvVIS5Kgq8II4mgpT/PJH09Y6FPRg8ycZvEdZXkaFvNX/m3yEi3ww
8K3NZZwgFJcFC3RNOG46uMnXmSGGqop+DAfVocCa0JP/pb/z1F7jgo+i0ZeMvp/hBKXXCPLjygh7
MN7z/HYZBpfrNxHNskskFDckBOH/V7w1alev9uIgf70bq93BJ8ur3aCelUCg0OLnvRFqbKC/tefR
QvFGUjXIacT8Nw6iP66Xi3myRVhNjQqj15JMvDERcVdkzf0iLmfzQr0ZwtK0bhmUEnNuuibLHEKb
gVseYu3BrDvS/0aEtvVpyQFA2vYHdt/5Zbnm+VRYB+xibwTksg+SzSEyi5QZ7gnvB0cgVgNkiXTD
HU38JU2ykRGrFokTH4R02ehay011RxpI266mVXziJk+j616aMeRpeZcOoVncmYtYcye7BC7tJYPA
tIPHJGSzlHwrfksrtiXIyULtd5cAYYU5DGYLRQyOz8t3GO3CqdLmQzUVBtCxAB6RU4PgmHMS54rd
v4TrB/fAIPZCfiEY58TNQO/YD1RS5M6yL6KCZMbGAVmWnmwbmIQSF6L5V/mdga6gRAjjkDMeNngH
coRcwP5P+pD3udijobbI7gEH91k8995d7+mMFB0vl3AeJg9uFQrw3rx6l2zLNfyxXFjCM4gzPCbt
9G+WRtp7oSEgs8M3VQbhHot0F3UsANk1jX2mc1w/+ECWP6w0oAjRXNS4/Tod2TDwTZDifZp6y87H
+8+DDSTszYfEf7/AYvGrZDHFC/bhJMKCbRKHiTI9ENyiTb3DlKB0nQZskMV1OAgXWErY9Xbe0Db3
/k2DyEOnIRlrrXUYBEDSVoE39nAKo0WovXhSEm5/64BcTX7LcoFk6Ruzj/7CL5zUQvJC1Qm/tWzL
snMsk6pJhgszJJ324zBBQdHy0cfnb9LCii9JhHB13cK0HOMvsLvKZvQ+jRoULdmKQrRLSgXPsF1T
fusL/ZpNIBxdgaiQVJgDSEbTAZrKuQYonYg2+m/Gu/H4qD7CaK/BQTEaBUzlrDH/n8Cw6bLVWa2s
3NsXsxsC4lWaCj9UrhSXyYdcqKFgoTQ3oI1FyHXdlBWISDDQMIJooNYFBQhnLuoHtbre76YTAWfk
wSsQwN6rABgrO9y4rbSN1AnEc/h4KC47Zt3UD0YNamMCMRIrpb0ofI/5daYbSyVxrhioeabGGZx1
DTRAA9oFWsqKOshQwQt7r5ZtPFkXy7OFtfCmEPnKJjCcz+Nus29V/RlmLqUHvt49EO5DdFSfshZ5
3tISPkfbYJETlGIWAIxSjQrIMncGxQ2WGwNTUOA8eRwa30orLI/S/7R4XNMiQH0HPCoFoXEuq5qy
qefokxBe/iiyG1OGheDl054mID/anS3EbxvyVq27SJQyrWf+Zuq23Ta4VNYBzBNXlZaSOsfgn1U/
Lx5N2yPfezl+EkL8PGrqWuE7kDFAJkhLJNOIJeRuiESXOuIzGPTVvGXBNG1kN0ueK9VqP9ts11TM
1XZ5FIdFhlIVbDyyL31ZltFHLOmHWDwH1c6kBZza/5o1D15cEh54sTpuVbarFmvrA/FXcxNLPjrZ
k/9M3KgWWomr2YpXlldzcLdL7Cvh3FvmD7TaS4Gy0KoV2nYTvcQE75qMoOMUOxuUSFhTLqCdT9wm
8Dmg2JsEDaKw0Tmy6VTlUD27zm4F17dg+klP0QD+wna9E8GwAvqOLu64EP7QUxb91U65eKlWQWq5
FQ9Y6B3kfULfcgMx1FS1ZRL2s96A0kvhJu20h0rA8XGILs1ytLHV5kG8NX6Rbtb55ERwc8n5VsVX
ii7syoyBOS681hoVXiq0fZLWNeD43Dpw2Tsv6WPK9MvDiYA84oTPjR089uDMgM3Hayy+V/liaO/d
WUixr3bidb9f3KQXUJ0JVfQm2pBHok4RsxISLlaznk3vWg9V4cb1pFS3eaZOJmMWMewNveMJwVwF
taMGlVOdDGANtK+DPtOkZWxpg9Rokx9HJtynVY0e+24sap37srzPiGSB26wNwBXBRM/55D6HIbNn
vWw3qJoIXH3BIEc3HN2Q5TdXdXXPaj4E1/eSCjOGX7IH/IfvxkPigRWxpGaULiMOZsRt+63iSr+l
FhB6oZhBiqUWnuKXZMWnldv/vVuzKcFzS+kptsaOxYOsE8vlo8a8DO3rMfixWCBPBW1LyQ8tOCYM
2GRG7fu8wk+U1bvZVc98+kqgBWejBOUwVHrflIaf6jW+HyWcpHVrYilIPN/QzuZlNnC5jgCrTQKo
WWCLBMFt6YwoyK/9qoA0MoDZc1zs8cTjs3f8VP1qcwCbPhu6pq1fCGUWGDNhveJqkWEVQbUidJvf
N6Y11LPNkxIFGpHsWSPYhda3V98HpAXaLDdN08tXFwU1xG2EWHuTD01MoGJoVkjauHVfiPkqEsQZ
7ftVcGeOHX8obRI/1b302wBGLqX7loYp7h6wYQnIDQZkYxOHwXBYA10r1TsMt8UVRXLiiVK+h/rp
05hWrpHTR8Xxu+5UyV0SOh/GBTbD9SCKE/RCD9QBywCAtAQitk3TMp3eGhgxyixaVAhw7rBQaUqw
9LuUXLX/Awa/a0innSI/fUu5nu5vtthVaG5F5dTx0adAYEt4yIosfXV7MYrTc1Q9KzZ6ECCW2fVJ
itj+JQX5hPEnbZjShVGwaE8xdfmpF3SuJUGa35+vfhpjhPVpPugcohDx868OPKZB4DDrJroF5rTc
DsLawNbiwlZgPDn9cFnzhvg0jhpEIhPEL3iArOVWXN88J0NG0RFPhchT6C+kCa8RZIVTV9P6Ns6R
sbICfMebN+9tNYfZt46a3z/tUmGxpZgXocKf7CGBI9aZ797I2bFQX9AE0lvGfjNcURgaOdcLelYz
gsKtgUsIDsfuZAYeiG2deZATA49bMj0/EcOhy1VtAM/uZ1GXuMNXQflG6bYPukECmu2wa5aisYaW
PdBipeMctQGY0GxIeaep5IgqwyE0qxQrFefvnJRr3GRBLvABJK9QfYWXk4uTrbfwvXFDb3uZQ2PV
bTOX3mWH5EIqlOQDZ5lzivy51fSlXyuOcNBmoDmDjQCii0SEOzSHndwJVuIw0Y5Xe1e1j3h210NW
4mS/T8Oyj30lCNjVvOJDJUcgj1aM48JZgmQ2sDsIppVwmZkrhrI1SGrmFLICyPGkz0I9dSrCDLQb
eDi3tQ8QKKWuhMp3zALlu+WFmBHHRhTIeZAP2Rkd64psUF5c+XM5w2mwG2JKkelxkKWQ/TTziS1n
aeKrc2S+wO4lgzugqFcITUdZ8Hlhz/Q6cbJXTCmg4PvprmFtnjvq4fugQZ67ehPtYDAWL3L+0GZs
goHLJg6dwXzobrMJczEfUK7/58HpNFGU/Zik6Y9rLV7H3ox0jo6IHcwzKpItkYKRa7IuHz7fIfxP
7kjptM25LzIwy6srI79YKI0Xthjq7g+c1o+/c2hGQogli8FDiJpzoe5Qg5YfR5d/6YkzOc1tWmXI
X++O9kyNapZBCy6OdUnqi8yNHyJ7SpvjyokYlYXw575ixAi0Nm9yrULT3S08sP/Mt6L4vghwnwZP
KmDXdsTIeyMespe531VH1SNMTBj3KmY1eVTv/6FDXik/ND7Iseg/LPKpQpT3qe/P0b/7GWK32LiV
+w6RXdkuo/HP10hrp/15Y8JVVOWsYinYnCShl8rh/nLVRB/Qw8O+Z/qxZY5Qrm4eovY8s7VW+Ool
9MeVcO1m9BTgD96Pdhs4NpI36u20u17JD1uMhKhZh4Xcn8BH/yEcNvsDnWc8XrdpEA6o0ULwzp2C
FspbYeTNQJLBuaJiBb03kqOUX0a1avsivIwDssKjW0W4uMpIZTf90ugbqbHc/3kI5Q6/ZQaDp/FP
4dXLtCMiek8sWDafBfY1p8yDfoLl5rDKLGoYDuKwFbe2WK1/OGoCGK3Jib1w8IayWwwxj38jz7ct
9Bv0mSTeO487EF01usB7Cl73GDd6L35mN4sBJktxdJWp93mPbnwEIDTTS3EQ3Ze3+WFM/zxNvWX7
6u9+KUFXlf0AIUQxtc8+tMMeYb18W8GVCSw5OWF5SxF5+APrVhdzatVCJcSi95sHEGFy+O3wu9yv
RyYZi0WQqxr0toDmYevRK/4SMS7ab58VmAJJSnupCDpp/a7GgvAGdS15PdtXqlgILI0uRSl2K30o
xRcbse/3ELq3PGmdkKeRuMVHKN3zK7jhCQRVemH1FepYkyQ7/RHFgNlfXAka2uVkw4dtxuvJF0yJ
BbdrYuGPj9bwBy6qjqsDYewWjet0B03qcwUz2ufWp3IAcZRplWL39pRHkdWl6dM3BuYc9A3SQgIh
KnFu4mdKXedY2Ly3FW7NI5amsAciEiqnNaokPrFC977Bf3iBxZId+K2Tzb+glpSjPkVPbA3mj/P3
Egw5+VEx4xVKY4sL9RjY2xwyIlmmcAYfRB888SwnksIEo60KIC986YmfieNuwXc5ICAUIszr3cNS
l9nhSybl8uF3UQUAff1AsIbvGQTx24dCEnxGCHQIqMtzjxKdUgikFA4F1Q9/sQrCVyVfm+k4rFq9
IUodCjqkeOI9YLI1UGNf3frKjru9bprNUUCA3ak42Iah6XiRythFEFNYiDQ/jT/nalgG1THF2fUR
06/9kaTPHlAs4Mn6RlcN1b6P96x/j5UyOq0NZ4cYHNCCLZGVc4X1BqbqS/yF7QzztQpZSBJA4H8s
4HqYQsPC1aNwLab0z+cfCOlkgGlFv/hBm4curophoXTo6w4BArLLv2JrBO1Cr0S+d5aNh94/0EX1
4+MRUNPRNZdBNqcQLq9m0Hv7xZSf7POZwIpTwLpicOX7Yyks5OsKOGR1DADeAhWXZxHYD4TYT1ST
Q2BJVNekhqY400JF1lWjI3t+SJjnCj8gcSDEyQKaphkPc+erwgHk3uI03YI1mOobI8YkLZUj38M1
0pUTM8bWZwmWyn0BvxljFlsY+X9SNt51YLKTf+KVancseLjb17P3uz8ktw6I9kXIYvzMhjpl8csY
JePOnuWu+S5BHFCQzsK5thZKhNNS7pRRfowNLmOFDT+oTsb3t+YNuceEG+CGdhoR0dAxhgfM0ll1
e9QYiOR7j/VWZQFKluYvYW3Add7mwYNkIv9EBgqjfFNN7+NRXvmjlTB72Ic28aZSonvJ7fdneHMj
yWMkyiPCoquzxA7Yvb3nAIu007bjIGIE6wQ3pqK8R4v90KeiiSdyzMecqevsNYIjibjm+FrEhHM+
7/ksgUVzZImpK+34z8laNgLs6QU9UbWINffWLDiuaazzK9ZoKNgmOqIP+WJJYpvUu4F52p1kSK0M
PRw740sdoWpFPSWFDEFEzTasBTTNK6xMm4s+F356ITOY5AJ8hWbg5/bHuaU97HaiClfMGqRc86QI
fUREZ8YM6qrubd9co4Hbq9FDe5nhqgizJdh/Y7OLYfE9ZKqHfA2NrSsiwiDua45LNSYZgV99j2Rb
+0vLswiuCOfZAdb9JSWXhpe3v0qFPXaYcwCVkKOMXEljnWa57gHtpd6Jsu8pFC2jRoA7BiaIVHBj
VL7Izi1MMiL90uxc6VB+SLxM1AunuVLKzpHsSs7ioqaXyhTl4I8xFe6eZFgGHXVBmPw1mjz+Rjwg
38ZUsmOuZZ9SUVPnWWmL6oi5VO9wbarHcsnPTXGFypSMQrG8yeJBwG8mLvPQ/Ue0Sjy2xhNewofN
iasQghqonPLSF8qB9UwCm3N7BNA3WpfO64tj3w0wFi8M+XdLEgCalW4lH47BPcEPUeXaGCwKw2hm
WJX4juw2iIf64uVGu0YMJreWIy126xnbsVz3HTmfoZbkYjNK/kL7y0swbvOz7wuk+77vHoWr1nHa
AVYV1V0hlEp7/Y+MquDZ0zRRE6KqUWEtpAmainpAYNo/UXRML/gTXXU7z5KaU6l3rd9PIcrB6xjS
im6TtFxmPkQb048tmd+ePgPldupxQVmUVEA61VmJAIq42MMEaqhvuTFDAh53K2K+yhTfKS5vadoO
ifqjKU54DNa7JqAZ+jfItJjFclVSNCyzCZE9yEGmOslk7kEWAOonG/qoMAGseYvpzsMoCLCkblTq
5dbrvpK53Qqc0+kjdcLY/ipfBiZPziW4n6oGZWfkon0azGYn8Ux3licQ5N+kmQjYBERQwkVvsKw3
TIZIbFo0fpye5Qwd9j82ToYAwo8Pd+50xTh0RE6OGHvJhkyWbJiAYjiUjzuBFw9qiwfEt7OsqRiF
HLAe1SZFrh8COI+9T7xfwpT0HhDIoPVicZdPzq7nC/hLW4ipfzmJtfHKD47VutztF6rAnNRrYrtP
nDOl9B1bqbplYnKtM6B4FRti594vfFtpcMhqwpbPywQuvqk/Z90CNiazMKw77lsZh6VRCznARLNh
RTqjaeURYrZAnojAQoknTzK680q7/WcnxMEYggF5GEgRm3rSmpUxTJIsekkbB9m4ZhlItKx/pPNK
Ciksrm9WYVdOIlW7//nw/6JawAQT5M3o8SoQWCeKPfCbC4c/2ttmHH6gbdzq211eDBCmn9C7W9UB
iszZqO02x3ybJnLld/bQ9TFjE3FP/1D4vynPFdSlnKavt0mwZxJhrR0cuABPtHwkOQpEESNgXa5c
MR4Vy4TnjfJGwNHyGmzOcuCnHrzVNhNbYE0itJo1Ce73UY+Thm8xP65GS9PQJTHSvNz1/fJhyXwN
ej2l6nz4uvr3a1a6C5GbqszbuNWqpwMjtqaLmBGBfyeSZyNLjObo8Dvp2V6YpPh14qX6+Njo6oZp
T02QoqObpy1fmrLroPwRW+s62JD/17eqYahL3qLfVSGoOpmn5nw/Mz9JO1veGldUtZtrnB7ZUa46
5Yub/pE8OeZZYyP/nColPSw0CwqWI6tggmC+SRVhMgXbppguQ8Iysu/4VEAJLM4KCm3Jk99zOLrv
31oRfg2ocTSTmYomGMpIdzr4jV5TSbYAADa45iKGVg4J8DxT7GioKZ3IPrRRAAriPE/ZWjVgAEvl
kfXS5cKBRYPJuthkBOC/zQUPPP0i+h3tFGJ7rX/GpvAoCPALpxC8tn7uvyQcliTxEqFRk8plfESl
CrLsx6xN6LlloAF1P6yOKQ/VqPXqRrBX0xOZucN1Rpgo59UPc8RgwhxwepMlPrtgXcz3iITM2Ica
Oyx1RkxVQsU50Xtsy/gMx+kDQKmO9UHL1IeHFzYo1nda7GWz2DpqY0bMHDfZETQqvcbdlzoTtiqd
/j1keQfFcsoB7wGwhVD4zDnnLKgF8O0C9nBKBHVzGgsi9xAYhxXIa7hVCY4OgpSXqk1zdSqwdK3n
LaNOy1GeOUsxsXGSOgU2+WIyL7VnDJT9/G/s/n4VIL4niV+REzDhxEHdu9gc4OeEUzCj55ZRUwE6
UiTn9cqNTbcmv+VWCF0r0v3YpLO4ITiZn3irOpFE17v8nb135Zxz9a95Kl40I3Od2oV3/zL279Ou
LgVcsXTlNgUPcsV+a+JThqKJOs0ZV98Y1NoQTV40hQ40tcTdgdMHskoY1FgiOWvR05oauTTz3MmI
M2UG1SbeHFwMfjfGS/lanFAAJ6taQr/ox2YetKfyysrzYfS/sVavE2txApcxgHOY05TNsPjmR7up
WWCmLF0MiWL2PFS7tGQvL2lBTLzHpPXaexykOqnTVWYVVrZWrngb4nTvbrsCaZTu3cPsXT830N6A
zhHVvlpchBnmqMyIYsoZfzEKvwsIo3LIro+5f6UeNB0vUNqIqgDpuvMLpe2A/5uc2fEhIdaAF4Lf
WDsy6gfn+sEgJzf4WEImHiSJNxBYwwp8EY2aFf1ZBO1eKLzx9yPOOoz6h8vJa32GYYluW4jMFxqw
vU70BjoeZe9rbG45RlQxy/X0h89TasQG9doZAOHDT4L+5fMJs6POD+xC3L3flvv+kKa7dbRmIXM/
R4Xgp96W01+gLfk7GoSb5DbphTEytNEhZrpwqh4wFgUIaRxzWQZhFClHPCyXfIjAEqPWGORFwm8v
oXw5qKBXnnVgVbhsR0sPycYdczTads9sFg5IqXfREDW6s2sKLsQj3Yxnr5Fm7hpHajw35lfctwjt
wZnCpm/ugfJvA2Gs7nc+HLBRaf/sIaZ1+i90y2qea7HZLvy8JWVfouADzUpzPN0oLg4L/rv6p7Mh
HBYiTCV7RjYDiVYZLHv195HoT3CfErDwujjdR5kQKDuPMx73Po/a6WYfSjjYyNjE3RRqb8aSvhwe
DZhPIwJRVvyJDjDQId1TCWe3Szip07Fj6pgc4KS36l4mBHSIJLBpmtr4Yp87fO7W1/lxfTY00DmJ
SvGb45qmDQPXDrsnzjXYkdfUkPBpsPbCAG8GDuI3Q8G2r0vOeCD4GUMyU3BWbgTtgAOYocmm1Qnr
iLFvGwEAtokiiB/+T5DEXHbK+0Mq9DL/ZisBNg+vtbXXoxEr90pI2azFmvsNINCdHXgKxT/gbY7O
4epPtiEZ9HQOArGiedyBWVW4cvQxL+lj99bu2uJQCEhBBDrsRwkzf0LUFpbtjaq3K0Fb3QpiEPEa
jjp0qatr1yC9uBLPxrwmQ7PmgNQ2yH8O7AZqoBAgAZcu816o/0ky2auOn40sA+NjcW/kRkzIiZLF
rx0RvIuiSeVjqhOPiyMqeClICstwYlKyR/h7xYaINI/8k3i12NRMpt+J7i8VQZfflCchhumytfHE
3mf7i/tpxdznbU8xfc8isauRkOHmnra5KfJA8VTwAgbGfBARbUqE14AkcMdomGOQ51sgtlSjM5Qq
2FpfRsEuzz6FwqEBXoRa9BMe0kwRhbKSO2EGHhEepmnRgWRgqFAEwnJLYf8O+t2FLLJ8roYUENYt
i7XZ/VyPcZ1Mwp31YT4Gs+qVUtzKZwhJgKQ8zxWtK6Z3scdLF7O2tuGE7eVMTYOPXoMcuiNCpBNa
7S1xRCRKvrabApjaoGM2xGdnSFsX6CDT9NLGglMSkmvBFCO1tdqyTMQtnqO84F/QgyvAe2F1lp62
HkQJhgYNg1w46Se4+f/6QQklYf71T+lF0/+Vn4nWaAmB5KODytcw/+sFyj8WDIhuRn3h8OglqOwd
/UBlgIzZOVZDl1NVoEZDwgD7hgQ0Um9AW1L+qNgvZj9Nczkri/ExSA4phu0ie1PWZJpeonkBwclD
gMGgXGno16z+IjB4+gRFc85cXV5HC1MZLJ71dQ54eOIHUR0ejLEJoc1SXvHqOi4InJWL0tZN+qqz
AfumjcgtG+2s9KmdGWr1NGqv1surcOnowSVAkO8QGBoiXKARcyMgB0BizgCPPnvN7X1RAb3u249H
phPw9rL1id6ce332rad3FVE6gw31nJp4CpnpxEf3oIProySeDmyVrr5jvbiL0/JC6S/KW9AydxRV
165ehCNowxVm9VxQdgt/BX0x1yz1bKDgjqy6Kz9QdyAiQ6JXxryBjOJLmh8epKm0FGl29dCeWZak
pxNcYRB16ZERRlN26Jb7bVkzn03uG/HKOw6s/F0FrrLs/A5Igpah0QTNonJdXk97s+1RBvIh5JQy
6U8LYuBYrbzBu9rghOqGO1CZVOzLPDZqVwn+4QRQzxAMlQc+3XWr4Df27aaPFkNYw7e6vU3mNajD
zTy4lAOI2Vp2/1JNh9dnAwihEFzP7cCPO3XrVdG10zYcYPx7XTWw1tPf3Cl8fwLKP14ZxuaukDw+
yAuoSqHyEkyAma6MXfpEiszVSB1HrMaHzkmtg6J0cSCnup9F/7OFRgBiyFGwNld/1S3WjVjzAEQo
qvY6OBPQ5ZzLBn3Bdz88VzghaFdQSWae9b6GCc5loQd8/WHMUNZXTgKpUJiZuP9MA+nNBCV9sFyW
xG4vNA8FFgym9Vk8PQ4b9dw7VexWeiUbjDMtZewS+sa5QdwGdEXk0xSbU0ZHFKzDN/CCpvw0oYpP
VLYOK8yYM77MP+4FAmpN5Kh0rwlxVt+npDOycEW6sa5Hb/8Ehb5fy6CyLPMG31wVkf2ar93vi1k8
mDNGpOowXrJrkJ03X+06qBxCHFhGb6NweSG+os0/vnV9PD4KDLDGr/WasAjDNCKkAqaymRAA/X1y
+Yb/TM0BQzK3ayyprL1DNHCN2psyqHwMjKXHO/XBkjqF4IDVsY2LeujHdnj0hAFth0uKJsyuvT8S
+qfKPp/LwxVAysX1fKgRpXwBYDZW0QC22Ro1aGUutEj3STAeT+uy9cReiNgDfyQplDgpEZL3O91e
gvi0xTyP8EGsm+0ysw0cZ9mq1An1nWgMRTjInkrbUV32plFQf3pB0OjHRGjXzOvuDz+MLZjLgE1q
VfcyNsqiSzRUt9nU1U/fhfYR9g4ZgQyrNJ3v2jY3ed+dwPevyn8IkYjn9KqDO0Wr9Z/jwPGaq/Ov
0pcVw+3OgGJBVeW/epS7ftxkrNsQP5VU4wcjrxXvf6JEtlBfxaY/mv9jzLy7CO2UyukxqRPsV52r
OUsL7BF/wCI9SFBNrraU90yf59BoDlUz5S1Id9wTS0K+zAi8JSj/N+0tJ3PAms9oqWw8ML72P0uc
hFVxbCM1XJVJQaagtxfCH4Es/KGCEBefQd682Oh+GARqpfMM68V8NkcjB0r/7NM51uzHxLVQTEgB
vtvkpsTnW/C6nzlwlAMiUXTnvQ4B17gBpZKBgLt6x4WRvBh4v+re4fngvcDU3A+bhn+qYqEauFZx
L8hP8tyKvCmXpNng22VjwW+La5e25L4DhgGY6AfF/mljQeKPAPaKcmJaMpd8NbkIexdjHEk5dOCR
8Ud6FnwO1pxmNW51eiwoYIyAA4ohNXv8oi89TyWNoI2cVDSHdrk9ov8OP6NRolBtrzyTd9wuJn9f
rsU9V1/oxWYELc9kKzjWeBUmsMTfndlc/omfcKa0eU9UrtwlSj2PPk2HQpvjlyLhMP1f4+KMU1zG
K60UgqshKtDBubHzCONsAmzNomElPyq5VJ6mA6lWEWuT6ShgKavXL2YHj9yfMFRXmq60JmP5wUbZ
9tF72siV3grJJviMEkNOublxKjHlzjLH089sPMNHnk/hNMQbRYEqCUjkDWjcp+MkfH3KpK6DbOm8
pZDRQfGfL4eJqfupJqFx5HPi1lR8uKESOSYqQtU2dyXwJxBM+m6SdBMEChm4X4WK2Mx08qcFWnhO
IMutLosc/xSgIKb6G4QKT5ZVmYGTuMejVRj4Biye3E0fPxcfBOJJdvy8M96fMNfbAZl/VECDWuUx
u/V7iIkUvF7WuOwudje4MfyDj+3eyCZWQctTE2bzAez2TzTctXmkD2M3DQUePC8p4xBIh7J+7KYb
cKZDPUl9/fpk9TIeq8uDmnC3Ma64xgcrHcAvVCkLPws6Wy2etNkcneEeMmlGRbJr28ww1QGIGbhz
z/6NzQrTGU+YNbDqdpERGZ/+aae5asMgPpHE/4s5vehRDvvF1Pmf+zFyfIDk/9CiGeZc+9QLY1v9
Dqm2VbUAwH59AsZhh5RXeROYMsdDNigCoJmKFLL1ZmnS5DsMqlOy/neU04QGIuVpLJyCa+N3DHX8
uY6/F3/9DPan1zoIar4bZq/7Zzs+G78KP9b3z/NQk0kZ4NDKMLnrOfHSM4I1rhtuCewAEw7QnPDb
b0lp0l6lC9CK+f+mTTKe3GQtJn6thUlFpGvgIcWeqgu6rZUmnX+PC8OQwqiGlTSqCCMgHW7swM1n
SEpCAnoHn1TfH8YiUZnHxdeN9Ui8EwBi+VVTJzEd0PlNdUHNdCY7b6hLDv/gN3BLng5a3IGpdcXj
Hbln0qKfgW0DLLBaTeVslh+tQ6RF0NjChxQYNTsePoK7R4DMBAItwmiyp7xrT1s/CUYjijwwUjzZ
A9qXSvJhsfnxY57wzz26QalRVtKlA9NHidBVVAJ8/fKdEuzgG9ZI6j6BzIoqsr5LfofB6uncsg18
AnfBlxPaCtM77XTMNAiRxjiBZWvvLUCNwjgXXZwrSlKt/dLNW2vuIciB1kA9QoTCTeWhr8l4I6Bp
wnvDgXNgPCG0sf7WNsh8aI0qm+vI41n5dcj/pLWdsaGM12XE0r7nYkSCltN0WUiEu2UatPkz3Mf8
4YvbDDe10s0oMQXwNBDAUBfMjEwjBWEQ4X/u4MIvk1lcuj2fwe/7QibaMiOuSOU0mT4huCdazO3N
qKjjCpaYkfSJExsl260vtPK+WOld3M8I9uXOjGz/liGk021gQ7llg/ckYzSAkgRl+EqVfIdYgs47
tFWG+VBtg7WJaSrHqKMB01N8oFASwZIdx/Kl5DHYYWPyub265z+a+9vWNEw54Y8x57Q5M3jpx0Rq
GLsycNiPT8phQ6q2C6a7okU7NFF2c5JO9DxGnnM5r/kcxSioguShdlEifZb1KbmnIfhmrqyYVLc3
TKaqrh3ZAEqn20BjO93E/cs/nvH/ofDyOnBo525tLxYgRZr8LEUMBKwUaBIv5u77a/Z9OT9Ln7ST
1KUFvAV92Xqb953dmjQG+J+7CTFowf1b4oENQ5WjdFQg4eG1g7/dbeXJ12H61/33sXH1I5JgHiXs
so/3rz5VRg9d7L4PLRVqv3ADUt4Vi9WBJNpPUS0oKByAz+98LHdwcIZG8m0WHzuYjlfFO1qe0Uux
xR2+F63kU6gV3sSe/jpeiGp2ahfZzdPpZ1ri1PG6kcpOYL0Eo7iacQ4kK1xGFp+pnwqdbYuinsr6
kgxE3LVyryUCmGJh2lzBi6monc7ryjGzexjTZvhUasKH1XqE44dxGr/aCK8S5Ctff3U8NOL4BwMW
IF1DY/6toTxvNcoAJQq8HgtCGDeDWtUXjdTJhnmoF6Ikav6WGF6qhBJTp4YP4nIVpElOv+5BEu/F
X2boP+CfsRP8EFJ062DV+89yPX6P0T1mGfUd0eBUK6WOyvex2apNX6ZSuLVHNOEN/6WAjIDVee96
IEOhW1Xihw6o1D2eD/h7dMry+Ac1T4rHmSWzN8WHkmp2uoBUZmW3nB26N+/ysLmX5WzafdB3UOTx
hit0qxxzoA0fsj0Py3XCIllJbWBCNM+4zPAmfAjZekjabaJ712rbPpcI52UA2yimmxvh+QtC3LmA
4M8Qe8E55PNWxQLjWA4oUBdCF5+YKXRlpAshfdTH9eaaPjfbuoGCaoaVCnuyRW7T56kttZEZvUUV
c660EZTQUStQXoIsMn4AumQRpLVIxhg/Uh6S4ZHN3izMQG+WL6DampEnWbHAW8i5r8UkeyXg5GMX
fOqRcC4RJDN3yEOPPfl9p0rTrj75+2Sn0DubDtTi45dmmg7wVtuaB3mAC0KqU0ywpTWxZCMqj6Tv
4TCo7q6Hja1dmAJHH1ywSJ4wAluuHmOQ8VF8wxiwIZDG8jL0fdHpxPQrFBFHJoTEDQRP2BTP4Zf/
u+6pP4U7KfqJ4g9i49zlchhzQ0wLQeXaeXmohgTIFfawsqghg3J3nSMUOUfFYaolfEBvlPsLbUbl
1fKDE23/MTDV/7hpeg5saNMawMp2NmHKBsgy9wAvwic5bnUjwbyPiho54Ob0pCdal+Zwq30Q+Ar7
I4pFx2uYo0kHStJ01YZk9K/feI67xbA/mJmVP6F7LHTekK57YCv28Rd8VdPoVPDMit8l/g9vnl5Z
Wj7ZLI3wF29e/0Go0bUL83r+hdu8YRz6hB/2DNH6eey20eNlHRodIAbqIiNcwQU9Gaq3TcHyUkRv
rKBw6ipxKFBBjy/o5xrze4fRMEqYSYGkmNg6MAyXbOd6p0wVMiag4bYfUw3IKhN7uCQcnraUyo3L
BJfWs+7rtZ/ayup8W9nvc3xyDTJh+wBzxEczPtVbVCxw8Dow+MK+P7dlQCH89B1XzIQlhJmLJrZb
tGb7xAlZuLqbrZtPCO6yH3UsxQqDFm8vxvRzrzBclqBXqSP85N5U2Uqr4R+fZ3LMev/FcyUO+42I
78QOO5t0uPoBr4Y+ZCjJ621l6N2xNHGz10lBBSSHZDw9LNA+100dNs4v+Wv2VN5awuVesDV7NyEb
F0g+WTEu0am6/x1Uafar+l3mQ/sYmQx+HsSWHjGM5V6iCYWPRTCqdJLk+c0bkVtNPKa+n4yrY0F1
60bcOlZb34btVZaZoP10avcWtBpeZm1fmGkYETe4ccn6oBBSr8OzKaJWD3E6BefinbJ5mLlmMbvh
TxIXpKdF8cJ05XgOFkVX3k8K5wD7fAXUTGPqv3MqiZNjxJQ8vIKxfEH3kEOl0IyvF3dw8N7kBOK5
r76WYYq0PHJzmcBSnWvZKoVlUpT6YlGMmhl4zwhN7btSdEeza5e9LHFGZeoao9Ff83Y8XIK7Vxhc
0uBxoLwG/lA+NUa4U4z83EKbotGjFam1+4YXKvrbaKzjK3r+v9BrBrwDJsjtzgB37sP262Xj3md7
KDKWmphnQPOPGOlA2IAvSUxcdah+T1eIsYcnF0jeZW/XQpDw1I/WrMpvuqDVQHFAY2AOZfPighIB
4LKV1y7PfgWBhSxm33BLVW9qnz4bqoWmqeDwMWMBiZfy8aBuiYghTCvRlV8/i00R/aGOXZ2WFDmX
25e6maGHCknMyvg7lNnBhZL2g6YbOyvOQVU6T+ctp64gbB02ZiQLqqhztIFCdcH3RulpQBgAg+d5
G1pU8DMhewG3pPw3klyGv+WdNKw0mIHylUgtCrl7eba9bHPMOdOCbE6vtqS8uAGWI7vjjiYmq5ve
Dr596G33uhJNb6XNUdjNXFcwiz2+bI/72HCmQDC8mYKHo72XUJq51mLwdqrC4m6rcIWP+EfZs/oG
yHKjUfi4dCXW1B5ZGu5V7pG5m6lx3sCYyok7mrWoS+XUpOrGQ1F/X1QS5R2AxKcHCTSlGjetFQb3
aG7sKPc8/hIuohhvofCdMgfxBMqPcIYsM1Lyx3YS4RHgI8N/Wi/O8WCta90RrBTMViGGQqI1j9DB
f03v1SFe7QprkYaz2qSAyFByJB7LwRITOutM7h0SBnxdzB78aF/zR9uE/SvnDTac5WYJXteFN31N
HDIM5g0On8h46qXMeiCVsewgP8D0+YCKERu0vjxS7/FcfZTMJ/+fgAUiKMx/b0dFrRbvzOCyVs6+
iWk0FFyNTcHoAwwYJQAuCdc6HlC4zUgI2drr6EKdv15skUzAYSqi40YtrmEXsTuuHiY7vvMeH34h
Smd+XHadbsMIaTpRTOX4R7LZ3mKNS1D7XZw8DEpx2+aMcU9XkzGvmMX8Qg+5cY4xQklMug2xBFLs
/f0R1nEIXggWGasRo/7FtMzUqUoxa4D1rbC0ko4WSh3oQqfVXWl2Lmf5ogO3P5kTDScyBBS4rVJK
Q64kf5BcC0mRERmcqFJS5E0W4LWanzqtRaH2uPM8Qbsye9OydM/9buz0Y9BrAzHJELfPw/YCxw3K
HL24Xazy/XD3CaYErif68oPowmrpFKSGKhpi98Cp5Z2v5MA08kDNZLofzPrdRTft2Fk8zgUZ4mLN
9NljZddAFqzzK4QAuskvTQ8njf3LBnz/F+ZnRwNwxqrz/tZYLQzmyqWHeuIMlHq7L9jC1bSf6oi3
F2LW/zuCKE0foG+ztp1rz0U+jtGSKTtyqTIFYKiW5c9SR4AtKlQnAetfjRx7p+9baxAFffDZxNDd
GBoWFTlqQDtyCM5qc/DtwNckMuqt6ovcXopupQsJYNW3quuH6wJAe/fRb7OVTkquTubZ0N2LRyxe
qz3s0xBOgD66ier02kz4WU7L7BSr0usVHMn2d2xXVcZJhzLNMOG36eqPdlatkw/f/zW1afBGRfs5
i779l3heBENiPET0Y7jHrdheyn1aHnI8HaSY2rl1bupp3Xya+/aER7cg0FJYWCbZW8G7w7JvQTgl
1eceUCU5Ere1ZghfD6OsYm1Lw1Uu9Mojh2D3oHiea9Lw+sY20/J+5nJYnOGVdd4SUUFWuUeSEEBH
Sif3K+kmcaWTmyTdN1w+UH+RMwVR9e+HWsDwWX59uFIePD1gv7Sc67oCgKG0HvLm+FgVkMaDyTmU
bBL+nsEItbuH26hs7/VN0hPnMWQOruWwxaf1R0Xz9Dy+WXbUjc8MBKYLtZXgvlibRjbmtkfIUs5b
eGGV+idOXvg2QIu3EeiFkXRqzLg3exiDSCVDzlKTzLNlQCjPvCPTnwes75lgrAl/ccITbSmkq0S8
EMQ4y/igFNe/oR9fONuzpA6WzU0P4/2/97jt7+EZgyDik8IOzef7y9QNLzAuvg0Jd/WZdmbCKezZ
cVHVKc8NEPH83fa95DgmQGvSesKddHQYftHwp+DBZcXRn4Bt0bUmAAyk7MiZf79xjupPOmlHPggb
ItgKesTXNBIphY3IhVT36R0WLDaY0CvJNDoi1pwYTqzlo2RhjT9o7dw2tG8CMQtfnD03SrCKbvGC
nG4uRGkOxMMt7BP71wGLz4IEdOk60EZAUaCk1s4whS/9FuWT7ilslEYjlRh3t16DEl7JJByYryZh
12MUkCRhZ6CdzTdgzYYiWyhbU7v/b+aVH4aAj3bAV8tB+hfJV2RAIIJ7OnhGGkc9heMAzzrG4fWN
kIrCHNku6YhoHqS601WA+5zF/yOxPKBSw3MN/xFWm89tJSlpdFKSbneicc2ofH+PF4njLcvivkbX
89WGpYZfwASeGyTjRZ1XHSBYWJgLIc3KB2MZ5gJAI+K1oWDMWiJRiqSGZdjkKxctfr+zTE5IM2e2
9WwfWne0UrJnqBl/3r0cwc2G8hpRrgWcaQX5JIL+1NU4ucK/3z6T1zJNzwG2bJldtz1Xa6QE4jRz
5Zp58OeSUU2m50pG0gf3dsm9vJsNuSKOyQ5sXGyW0hN+rnWPXvj/5UHvGpFJ+sidMt1gj8sjMpgF
h1pycfFEBjLjelyI5GvGCdY2Mr4GZdcnM8qOAMRjTXmce4uxVEoTVkcygEYocFnsZE9nJIt5BGIS
H12p3WqAiJcFcuibD8KknfD0qQyHEMX13JAbFE1w2m56cQJrT6xYrQsuBfvUMqIRsM+9dN5cgBp4
69qbrGXRwJ/moQNvaLLlF+8v+BlyO3vLjAv0EVMlwDJYWJ/lM3ZZI+8mO3UAW3r2aEVOJNnkr8uB
L3RaC8mV1w1q4GqieKPTwDzBuMHk/iaL2CD6uRAeFrcv1SMUqXjwCGvuUuNaggUkKPklGhJwlbey
PQG7Mx8hIVcsDfqhGlcX+dAT7Vn0sG6B6cIQGertS9Cs8+tEhzQ1rfGTuiIbVJQJSRd7diw8Wm7O
+y8SV5akcCojzrxINmVOMePPfDbX1rqt6zol7mDVhGWA5uflRgpyLyCDSBLMWaEXNfDzhfSU0lDD
iY3VguvNBzftUWAZZLhpBCpgIMil61ME2Gr41oaq7u7O7iDeGhOacQlKBNA0BbAnmfIs8/8gmUZ1
20rm0yu9MrKGl+JsAkBVxCwUS5tWORHkmY73RMb/PCZuv6ebhZxZ+dBZwBGDmJ8DyeCe50K+Ppie
OoELpV5LO/inB64ud6gnbzKJktMYitcEoHndCS0AOE2X+bNypFeio6pXKJ26+5q0f0NLhtfODvm7
d2D+4KuMGnerg7C8QqgWsu4metxwA+T1CrXTu//ZBzrlVrZ2H5UQZsNVFmSqNW5fD++yU6sBGACi
TRYdD5Rj4LZhGK3mKhz3aLxllNbcCwFmzoLfOlBg5quFy3TEorgfUFRfOfHVJQDNZQo15qvN+hyt
DHvIRT+ye/qS6EP1V2iGGInaildTYEnSqiaT2JdWGKc3e5aOcEhyIlWgoZK2CrRDiTUIR2qRp0oC
QiyvNGAYqbCn4MBboQL19aMR76C0PxL94Z8coatO3qw2rmbMLYdKxaKIiycWQOMJARoBTXWY/qgM
RYMXt9zk9ZB0hbnn8o+pIoABLQ7LJ2VG88ASryld5PhglJAWAErMe3Ek6hrGeuNE67QgTHmzecR1
pvceiHCwkJnYMEbpTD/fxKz7TQfUZIOo2J4cY6WV4us+/Qkv6iFIreZLQxC8pMjXz6EKqZoc7Dv5
PFAS6p8HL8M3RJYOuHFLwi5plluIfNyIEG4XV8DOo5eEwkzx92jsTzKaiKyfqKN+fjXMFZYszmZk
QIv1dQJBKaECm3tU3KYL7u5nSfkVsgmSyWUNi7lhnpmANKcqKLe8NXa5ebMQYEYjQ26PG4xh2AEL
ihemXvxpsGvtslRlvS1hGKDMxdYL48rFm6N2Ddr4sSJftDjJRJ+c3PBPuh/YdOyXfGFXQeT5t7IW
9/mQm1TFL3ITDdbWlRQZr3YIqeaJN5DGAaaARkJs0V9kfwGyYkmwaK3ZytBMuHN62SOmrjZa3Mwc
BtFpvgZmohJW7+g2w7HOCOe9kPnZNpOQ3CPfknQlVZ8x5rBmhppSb4f6lo4j5HLp7syLcz6uLZIZ
gjHRJCHFMwjqa0BWYIOLuVpma384My2LQ3NnFOf35Wzt030HDXfc59xyTZJ5tGbVvIEVWRmB5jCT
Ikv4MAfTWuGLGuqpy5v1GXbxFAtmoiMwHh9lkmRBIplOTJ0u5QkEQnEM5F5yxjF5k+iIXiHu/l1Q
xyb3Og9MOzK2WYRz0DFrOa5Oq8hkadWjFsXu+NvKkWzQESXMfH7qPLrmPoarLz/zLOALeSumLl1D
sKhwJprZ6GBYrPZK9+Et0/yjwDkhDq4iwm0dRZWaLjvBru397dIfXd/E3xnN+9VlUFGYe8Lhens8
Ma+oJ3jFYWGva5SQYw6s4CFdTSCssODqvBozOD0vFvHtQvJLIOD+ZThHTnM5v1caDEHjq8muo5Le
+yLWimXUQJkfPPLWMbQ6HQZiMxXwDigrGvIjiZQfTG3jQ75+tZ+VLprqC5dHWZ3vEjPT3gqW5sHs
5RVmkk44NCC9tBrFP47TujwILyip+VV7WwEp4Ml5E0jucnACM8kcG/L40hN5ku8Lsx5LeJEJ+UfJ
6A9R1u1j66zKiztfjEeZ/cj2CUObAKoO9X0LrHDNfnQ5mYeoQ6oLz3QAA02tcrR7X5jCov3ljnXG
asNL2rswlurezIZdhoRCplbwaHb8B27RVIfU3NYsQusb3HM9Ea/bZBoKEKkEFrJlNi1oZ1A3/9QY
R9e6l/yrJf44ikUTmiNYILCREcl9oyRUwzbXwNJC7dexZ2ZElHQBmi8Xn8w+aTkoeRvBkP0v9Z5k
HYlQJOqFt1uiZBRl3+L+PWov7gx6qbQ7bOB/OWG/8Q9ZLHmF+YY5xQwhF2iN5c+R3Voad/u5AKZP
5ep2FlHIO2Z+YUKhj4Kjl5IHdo/wscwRBZwGCmn5ZfNAjpK8eCMz6LPxqWRL0fuzkxGxCDMSw22M
Vh5JymsGz75yZh3arDWhf+NIWncfWaFNXpSFbWmFRUmkURPPgY1LXmCTFM7cdKFFA1fa9uDRcSCO
W9tVk3uRwlthmRUKNdPROCWRAJikT+HHgrYbFJanDqNwFnuzYAJS6SBJv60MJnmWC36JF4ZXpqaz
kzzwzO4p4A0FLCjbV8f+gkjAJf0X0pJn7PTw7tBa95sKNH1v6akeDwWk8iLre5ODzSgvfu8/OzF6
KdO2gjsrQunt3At5wEaWSKrLRriP7HGbmuNVX4coVGEsfagDGUnbCC7fplF/51jO24NLx6FYSJw+
jQx0hj9nn8ZtVf9+kxef0AyfbhjeTX2Tq4Za3JoCE4kRIgYzrqOaBa+VI76PbQEQTeCtlHamjNAo
MNpdgVuVrAgN8+HtTTe/W2mswaRfzeoU4DuyLMKBAP41bJqpd/ZMLwf/kNGpqXKIfJWlxt0hvHt6
siGbbl4JYGu473+QRFlSF4Cy/p+6yMBPdXWqXPYWToJ0J35eSQMgG3U+ZmVY/xjjg693gbzGajVh
u+qaEqHyIhcfFkPPCG176sYOpx3Ee9GQsI9WzNXdeV2K1Lg2/Vyck7TsFE1ylsOu2GmOts+KOTOq
3D5zxOQGaSLaqpe7vdcILMIMk0zsv1xqH7LcXxDm5ph8OWZ0k6lechBVYK7PI0qNgmB+xZVZK7cd
mRNacFkl+nokGxou1LxVDbG9qKBT2usa4YAdbtO3ZJg3qZMEJquGADi2IPfj3ru6r2ui/LcfJ706
QmT9L0VYWa6spYY7B+wX4HEp7gxYH7iH6NLOTKc5e7TLkE1gs4ZYZmvekgmMAF1JkN/IQ5vk9enZ
Skna08X1m7Ba9kH8XJrj2BbUGJ3Ph7/7BNT+CqrNAAmrpdpBOmGPTEIiArF/yhWQYnlwjxoPhkt2
16mgw+14RSqQW1jK9WeF2XEdJe8cHatcPDC4EM08qH23Da8xpmYXpFtm3n/gHShYmlKSLONZxUHy
ZhxcS9D2ghNFO6vZBlDG6jRypuZFGMR+bPR1zq0YO/4AM1MjTMZm1rcoBCatw2qeoJ8Zq7ffuV9h
27BbwzbLTu1bQhepa+2F57Rg6GgKByq+iDhhma3eQOEfBM7N6XJrOxTpCIK5NAyDrkeRFXPj8Z5C
OgIja9aivcGzSI4P9xR2qH/zGQbp+lOBiNLAdq96v+MMSRBtaHVufzNtV7OjsNya0V54hHMi7tGF
7Cv9hMSFQqNYRFXecOFva41LGh+comn16g46I6MBwIgPqrUICmXBS2jGqKJ43AHD+95vQagZCMFq
FdxHuPYZt9t4Xc5xlyqYwg/arZFVfp7LxnXEvA1YwNoim0Dk+w8wzZq+1ySNkdBps8YHxuEArelu
9XboXdl4chg2z0UJAfQH+AdeJoJj3eC1VPLmNJ4AmI/i78K1+urG920aa9XvzunR/BmABYAtZHEa
Yxl0SCx+RzLxie998A6kkZ8T3y3jjpTkdS55tUIv8Z1n/+/OfNYkd9OSfNJ0h3kMxv0mYxmV68t9
kSgj0/qY7YRwbdF9Kcqh1l11rmWev3aLTEp9Cg1CoZfOqqV1kRemes+sL6/7ZS0Y0VZENjvFR1cO
t9KBdprt9UmiwqBnhuoVerbMsId5mcCZytDB52Elbr6live+RwW9E8ha3IgdS4X06cJZbWyaztkQ
ZL25iMDyGxR+rGZ7CMrG/fxw72eJk7EvqGFOI52ie+YYAchc5M+1ouT5LqZMcQ93MEkxX/Nt2QVt
5yH+JqFnYfLGFAviux1q7miVir7zxK6WWtAa6GZtTNN8bzSF7tXCtgZeMJWRe6T/tYlYmOP3/yjW
uR9F7QfpGPndl8WZpqXwz/orwSHUQVuJXpdJkAEaTtKVx66mkmqRTw/69gvuLnJdiYc7CVZYv/K0
tiGTaocyu9oFls4vrm2f82lh2lQ7svhRMQxgamgVhwP+3Ha78tdL+iggVWBPm7L64kY93ud3DuaL
r7lnp4gECHkapTKcQZtgcI7io0/0vkEppZ7TbdTDUXQlKfnfWhRrmRVs0M4HZ2NGXVs0zkWY4VmE
7phP9+FtnFsCdSMTPODP1Z33uGpvHoL0H+lxKLX2Y5IWh8DbZlPrXA8LZzyHK0Ef82XLTDo2KyfA
DhaupvVhAL0V8t6HMStyraei/GJESsJjp0nxMr9XnFGMCmNeNt8ZbX83R5buZYvxPlYpsgmpaYIS
GnfS9IzxkYWgUSZS4aJqfu/77Ei752zMUV1V6OaS629/qdY1GsBVc88fZtRgJtJSRUnxmDKdNKRz
Pv3AtJiwVZAcZCSgxB+OquHXqWPy3jOHsnbFSDCXSMLFPqz4D6EWuNdrHiVpCh2NcIuYbUFO81z3
8uVTloR98i4vHXFZLe7r9SyEZUL1IYSVj2tuo/JikcQv4jAE0mULAsxxEDbFWKgnMHQBK/LqHShu
/X3ypI5OBD26D7SA5roWc6D+Fg7EoeZFso73alhUHWHs4NS+zYO7G9SqY9gfAaBhCy9sPdLFqIAD
duP3yvEArV11flvlFWaZhGO4BQHO9ah7b3nRvbYHw3+W926cyq+SioMlhkP1aeRXRUpyPm4MfSuE
tNZ2Y+VFnBRbPyvTIHOXP4hZuUz9kjB/QD37uMK271cgCAx2abcrF58OuZq8BCfIPu9cAyIj3HIH
NQGvkaRBOCZxwO7QX3sqBxuBeQOs78iAov9K7NosmqS0rFrIKcg2OJLNFXdzsx/T7XSjEV5mviYw
Cj71V/zb9v8aAFPWW5KIB/MYAsjNYtqIF1jvoanSfT3q7JJDArgVsRQf5cqjQl5KKqmCoGgqJXiY
Q1k8uMs8U+6LSrGCrORJXhRj2H3sS8mLAXAuR2QIc41816/0htxLNvWr9Mt7NQD2dHW/Zzuj0Gxz
bkB+h+FvI4udIkV4ImhoW+FRgn86koRWOmB+TLUiV+9rpRGHPH4YVRdm19lseiTs7aYHwry0ysh1
ejwZ00RJOV+d/FqviYmucgj8aFIatFK8Lx3X3htSyRc9umDFtoJL44RueLNgFtPn8dlh+JnEzXT1
QA3jCqpdlXgqEpey5VCRjXcGvGf2auOrg0okziFFiv5bH6aVlcSzdaN19lbolJiGE3Oimc5TbP4h
xXVmC8CoKB2OZIJhB+q7gRBphBVv+VEUUi0rlqFV5Iwjq9qR3E/G3+ds1QIdxUXPaLO/qdkLZTMr
YIVcn+NnZXcmFd6QYkEP9QKlcqwXfo6hulLQSweJLKNqWfSouPku+egdBfRonu7Gp1OSb+z1zUmD
kZr5y6k8vQJ1leepy31BezhzeV7/qfpeppvv7CW/7arKXcTCjYVYLcFdK9382x9+GSw6TrY0uGWX
6Z2vJFnFu59VK3/ggWleDpxtlfhg3p59o5pHLeYk2J3CAIT61UDGpiuo4quANUMjS+NsbNs3DnkX
gccNPnW6Xt36lv0O4yqJ95g8peVcIbHL8spyf3/9Id5UYrKVzO+YpalTE9Yq/k3ORk6NIfYj80DJ
TtcG/Sh/boFaPKHPnVhd81sUp92vCNB8ZF2lNXPXlpLw28b65T0DeSbFu4iL5gveimP78WgBF4Eu
PobudViYt5U=
`protect end_protected
