module square (
	
);

endmodule

//https://timetoexplore.net/blog/arty-fpga-vga-verilog-01