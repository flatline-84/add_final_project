
module hdmi_adc (

);

endmodule;