-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bBnwBVDcYk0Zt3l3dZ8Ibo22nfvTyXTN7m1c0ZLh03pXiSb0DKwzqLyD8oXpRMs3sl6kQjvJAwty
rC2hxkTdZ6NuiS54VOWIqg3xF510HrzHxiAbSSNaMZXgvwdmAtwwg3Mv8joSlS1UDHCL8dqEQN4g
3tY1DeIoA5KUmY1Y/BUtY/1Wb4/FmTBmcchBr3WxmwoXhlvtsmlXfpFQ2TWyUfJssB6VFaFeV+SA
EzQ61jYi64IsdWliamtMrd1CbbxGWriuzKnEIn3DeeRTQKo9SqG0B3RkFfyb7sJuL88VPue7pOk2
uqSvQ/fpGTVkChletBBrG+RZyhQuxpRn5R1A4g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25264)
`protect data_block
+1Gj1Xyrh0BBztAytrRgU4zGQIlWEzbkumfB44RS9B2+QToDiN2JSo0ELQk7F/8bLF58k/ZD3W62
+Mc1jIsZ/ZGpZWMcsnTgHofbRfDbT+6jSbulYAVzLlXlL+sbjVQAxnI8d0Z8e2LXCIbTsVJTt7Hc
Q2t9V62siv77ueS/QnH4XlsUYbXwjQG1QXWZf2fSuQZXxq/Gcr5N101pm84YtIgyHP/JLE5mtKa6
N4ru9h39GotuY4JCWMDwpcJl2ze97kiy1A4pvASXoUkq9hZsplMm8UpLW2a7bOXcgO+46mNPOsWB
dnCZR03Igiq9/wK19WyITLGQ8s6RfPYysWniryul2iJOItj7cdL4OhpThWsCNwIw8ZcOL2WLdofS
X8V+dLOVU0CXAy6e4zfmurSe4G4qwFtaWM4hIau5yLXeIo4BaCO0DPEZtP/kkAb25deo8Rbgz4+/
Z3PaU9qWCKgVo+nWkC7mllLmNPnJssz0SePFC3qEtRJyfx5utwYAuCviMK4MTiHLR7naXlu4MD0+
5fiPtGpgNUZUJCtUeFhEnIAxpIezZiK1Ujcxik/9MJebC3uUOdbIKpCpDYhUxQeZKQ0bEUyJGDCE
ds9Q1H0R9VUYuJlzAqufl0foI8vF1CoNRdlR0xw+7W/F4vsXXhXo2T0upEDmszoiJgguwz1tDlez
YYdca4bUR3LT+eTFIkAXX4g9W5deDnq5HkuJT4vi9/ac74Ovcv0Ojd9GGMR6Mic7KVv1uvf9cvkm
FM5vPnSZpfStnZR2k+Jtkn2j0snUGRcHTmYMOs2EBjhdpNt66db+EHQKRTQpIj2+CSCIGx9bEk3B
JrStW7XDxLZO1/MM4OBrCy/D722cOJaL8BIOxOr4TiqM3Wo+hbozfVBvcU5zoP769WELVd6pBX4u
F2Tw8n2UWaDSDYSxj05rvJQvoVtuhI1I9AttKPqE4RVjV06C90MZ72gfryMkYmpNTNah9EhIiUXF
AY9ryZnqlXfdqXApQidwzAsbr+41Q41uURgEOUIRWN4zVdGZg3LWDMHpAbI3/XanRIILE7e0Rgbk
n4TleEl8RrOiFqY2YcUeAE6hiR1BS28/PzDI3JoB/DmYdR1ocAM/eJjpdCb5Ts307YLvwXqZsjMk
3OicEA3lOyjNtmYBa3Wl0nO43mQ8BHz/CEw5jJpS3UUVrvhpOnZEOKY5kZANP1zlJ9UZqpt0tNhW
bnfMPfFVGYneZe71Udvit0evbrANnJwVlfcY0JriP1PnYEqnzHMOQuNQjPgfGSJhwkrHquK/QbYT
eTEzFwEl8wkkhES5woAFgK7EuX3KugZQtJYWTHTQtUf6GvAYckrYT5SmjdY9ZdRF6De/+9+6SxUN
t4q+AlQMGkhgrSZxvQ2HgvYnUIPoZDPoYq7zLlLcoD2CD1MESvsUwlFp7pZYanVabCiBujc9St0q
tc6gWIAuHuxW7aMXhE7tlN84xwZPF+MUBld28ptzGU8+Jln8rIwlwq0d065mq2y2qYyB2GR+fAwd
Nlxx23NYKFW1UwSnTjTxm+6B/OtiHWZcW9qYJ56t1U+EYHMh3BkRu4NEAj9ANuPxU0uVaf/k67B9
z/dXt35M6/tSCb/3MBH0RrknopiWUSelWGP1bRiysTdnopGK3QlZ6h7rNmpHobjiC3NAvDcrR9Fq
CQkjMmYIejD8cJNXU8uHFKgTt+d/Kdl1F2X/HVJHk7YqVofYbVbaHy65Ktllb4HzuY67pabV0IRc
Lj8z8BBauw/+bs7H+UtrlAIgUJV097waccRzp1FLvKAUjQWFZsZj0I8gS1tWFSfcNw2kMNJu2B3o
+k0F9IvGJfk8TN7x6eE1VbenzGl3wgox8HGvm+qB9e+4eBy79KPDAXbK/b+wWY9cw84cvrFlX1YI
cqKUDl0kiBMo2TEflPULuOlsQSvC+XGt4P52YrC5zd8T9X8b0qLn8TwHcl7voJ5AkO97SC6axO4A
sTmqwLPwnqFI/NUOtFpinhitDZXe0rtlOYNNr8NF/KcBV6YGYpLhU+7fKudkJxs4zo/uzP1jLGmA
m+o2zOaOdQhsibfJYfXclqnbiY0FPuBIOpMdfD2jHoph8+D/37ZHmFB3mRo+kM7688xaIA3zrvl1
0d87QcDD1eLIfuZOuaksF7yTyHy1ivCdQ4fn8k+dJtDfCxr/TaxSCZA5VthQV2ZE9XF3FOtFUmED
Xqjub/hFf/oQ5vbV+V5uaYHoIaOC7UZxlWBIP9+GPOgCOXumX2ntz9o0FcW375ac4ewuqcSBFDOF
EMukqvsBXGVMRoof8n2Q05ejjNwG6exUIxniPWMOeNZYyivtaZR84lbLUBaQ2dYmFsxPLsVaItKV
mYI3AvpCel9PeNxqNElCLbSPqfPHP8CSHkVXvCyA1gvcD8AJE1rROAMJIQxhdRC8eJYUg9lTmL/s
8WnFJCQY/JBrQYxQdFIVEQ/kmVkyXBHSM4QsWZrwrW54LaQD9VQ7vO5mW58u95wZhEluZGAL7OXl
PIUxsvkq/uyIVxlvcoHlnT0O9lBevhDDWSdS9nCu6eX3lMNWmNJ2KyFoI0ffCP+9uIp7eCMXDaBg
fGb8DrQCEtHyB+AX1nFcscrKhAPlDmQSOZYVWyJCCXsmCne728bhjk3LJ/uWByM8I+U4HEv/qGj1
HEiBQ4J2ehCYbekfWqWYKPiGE80DfFnT+pIuUm7rA4dBnw6gqCkP5dMCw2dO91YM79Yolyv0u61+
LxMVBAOj90/ZfvQ2tKzdVK2bxFhppQRavNzzsCuDhl0OyaKbO4JA5wAvA3u2eB8Ko2jm88TCLcu9
i87Ipy+8tY1wYvkjabSPQnQr5GMP1k4epqSjQ98sCDKsLsY3GOv6uon7jLmhHCBjUwlVlGBODo9w
2/Ka9+b0ZymXpv82RjEbbUfo/2w4UYApSPt6C/e/dYcmSVpikgjBOtC70G+o7CY0jF0iA7/agP06
x3OEOGtqFkW+aIbBAXsLZEzyOZsAhmTlApPn8ctAEDaNYu52w2wNtNn9bH+YdGz0UWY/RCU2hUsC
qTud/NfUvkfZtMOmGdSJ+mLMoHEEPD4CLFBmrrKm5NQEOUpg1xmdjehV77b0N3snz7U6FoaoFda1
+eGt803kX30fzmv9xC/weh5JvkRipjIqnlnVoNYdhPvzdkN9MLeysPTlUylI2Wh0CjJcUuCf0JiZ
1vF+kSExRAlXLTfBuyMNLGooo0IHPyG/Ho0qh18rJC8B7UusMPukPISZjq6om/z3nf01wq0Zvhe9
nevDpMxsaiCLOqzizQos1jaNgSrBFkWTN5tRXE/0GPy0RDPUSbaM8upKzquo4epmHAImLFYIkYT1
4wWNBSAgR53pdYGR7sDE5J6jYPzycgCRaDeRG42LyhEi7DMlQmn2Oak4h6+d9h3S3ePc+owojhqY
V+UVWK6W/cmeBAhjyVXKh4t4GjOs3sY6NtPZV9UJHKVk9g8xV1gg1xqN69Fov6Hbname04L6Ko44
OFjVqXxbXxQAgKPh9VicjtyeAXe6mf4W193TRFnICUDXvEWDis5zo+nFQA7AsUNd4yy0BLI6GYBI
HMygkLE/dybET0+TjYseAKSt/KIQpAdS7xdAmmApIvKIVse3zJEELXAOEtvN/PjKOboFLGomPzQa
+dGkCcBovmT5uUeu3XtEF5twAqofFs10s/1XiJruo6shGPFIoZDv8G9E2bb/qOtfNqHQfK0eNRS1
nxPCZJbXAuyhxAlNS/SXDnQAf+CUZokOoh1b/I//mWobFgErDFiECxxKQwiqADrxOYNgGv4FZl6T
yKybWzPMw83hRPZN0MozeNW29ict3EHXFeU+OR5FOdNOQWTSUZ+7iwQ+NcANe/hEsEJr7i85kstc
rH6TQrJ0ptxnXdW5PQ+Y8th4IHKJIGYZz6Thp8PxeoFoLLRyEWl5jv/hC1dicV5HnHvHxbI1MhV8
gQXpHS4ZM80KKjEjNLg1DwgnbN/h43jI+ZqEJ2sjuyOfX1JoIplirlRNZgL8/GcUqS1tVHK6Hzbf
4WUPLn3PnmExmAfUsyQYqruv+oAi6Z9A0fjrilqFJeL8ixkndhj5KS2Ru+BH+/NoMc6FG07A4kf5
8rNG3xxmltPVLZkke3/41vWbyof5jmJ77nf4PyXs1wLZjqogG5uDzWyOL1wjFeANPi9rZWLNd14Y
ReecN5juwXerJvmMrefX9HbifNISpCjKe6h+uTB7b9HOfhDj8bNneoIEt2cnjEhG7awWeuC+Qmfj
l4SJf2VOoa/iaBPw4YBK+ZdUOtt1GTvJLafSr82OXSwZRO+fcB+VLAdnvZNHKuXd9GvM3wae7SEt
7adPwZ+Vc0R7GcilbuUFs3fSCXZippevuwh3+W5aoTg1F/liftwCDh013u9+Bw+ZBYTFio7DxHsL
7l9BGoENuQIvoK7ya9U/VlPGT1oBtIMZS2aw3HPkl+rHGFGeJFFcbb4gDCi5n03jWbuf0ZqqrcCm
L28ezpQCXkThTvB5CMF18EX2jefl4jyFDJkQH0jrF1+vlT6rkk1Zr4MKo7Sh3r1psDoTPo6rN1+r
bmcXJBMNj7R0FsNREdwXXJPYMC5fx1XQqsMNGh8E/jplP8JeF35pwFjplvRC3kSINmfHFSTYQ23w
PxA/Zvs1bAmaEe70CjXfGnr2aCHQqKdYCjsM5+vHr4SjSP5XyZJrnrmpf5SbQSu72eLl7JK4szeK
xZ0mEMW+HiANtk5ojSV01/QBxBh/LpAT8Za364F+3WV0YWUduBwvxLtT96YUOFc0Q8CB5L9kumvS
kQei5wEe4Ayqyc+LfMOhI1bXoH4J5SEdgjs5DuEYEnHgkP+gVawMSJt8WuATGm14lum1bt8mSTOJ
r7gIYcYRwx9VKQv1R5/OfaWbFR0AsJeRh8SkmJY9oPoaK1FUQz2yxybLeJPiF7h/1cRfe9ZCJTow
yZ+gPe7ZeLENdePwWUs3tTPiRbHtmeIIV6zkBry3/fBl/fxdhOjgOhSwU8PuwVbP1CiKY6tWTxTf
TUrCsNdEVm2dfkeKI5DX8PdIXuUKsixa3lpNFMtGbV0hKrzAfxfvkdKAPriMINQfZsjdB8lqjmoD
XXS1CD/LQNjPebkTWhSR0rXntmmWGOuRbe7PYAzlvMVyQDJ3K5sya9QXHcrMliIMJDf6ZRuQGjZQ
1bF+tT4YwEfmBOwRgF5EeD0oNLX3jzUq1rOtLk1ZTsvDgM8IXn9pbz+uRP2Ajbc7rQ4ys7Kr8mqu
29VbPvmwKQmE2mQYSADXEtPSTpv1zl9AFoCSZVdhHNi2cuDwQsfctJx45+dymYvpDCKAFc2XGTKF
kMOrnsu8QDnXsaxnaplkJ9iNHsWTUgF/eksh0DuxCaKL8QE5J85JLWk+usIGVhLxYSc5I9FVpVSa
7zTA3hljOAv/dHNEE5lrs0eH1sYNZ4ne4uBvJ2Ms0EUBP4BASmKWvZPw6yC+BMfkBNX5wkhThUOD
aLDz2f2ujZAfoCpygeck+hX3GtP3jw79yQytk8kXcXISatgGLC4oaRvGWggp5jYuAxbQqCkRJwjb
u6rw5BuxuPU+B9PJPm7hG3I5libJ0XnLFLGQ8eCUwdUO2wKWf8AcQ4RRroQo5njajzCMxayM8q+l
XAHPw2mNI9t1OYhOcVp58EGAE3zMSa5iaLSDcR/+rtiEpn0AARySV9MhGD9OUfMOqsBy7fa2Mimn
fS2e1y00J9gHUoq7hUu4lJgQ5ahsM+LB+XyELZ7RVjB5hvY2QoWB1MHu3JwiFSh2PYU+bnObG8SO
e+GXWeWCU6BPLgOnBq7HupZKKCD8ISq2+1cPRysQEAOooOpLVupPI0JI05P0nTsFlKBRgn5L1coa
YL6Y9NsyS6bV/XfS9drUwdQaE5+kZFmmpPeH81xMoDliRyvHoEWOQ1weNu1+Jxd1w7WcKjIIvC6Q
s+vYfmqxiV45/NAvYKz4W5eWqIL8r8i7XuuipOcYzUAEcXNgjsDrlgmRECR2IfShyUuwGiPIMA7a
LqEtfFHOVHLaVa5dEhvNGDXYShwGpz5Q1GjZ29vGJbE+IEpKmVd+P1S8UhGAImqGxLZcIfK1djb2
vswV7fD7AUKqnHtLySdnCGxhAdql+Ouraz38SijYPrXnDKXQ5X4wu3sHSRhH1wWws/4V6tkFWkiq
m2+uNaNjU+2fIqIs1UpEJPPblr2eaOk4xAsasiZJoU3ZLoF04qZkK13EY/vFGe78ucQ91pPqaWtJ
ArcYoMxlzi5r8uceNQYScZyE9lNg/NGQii/CgpgvbpwU4GEUm1+RP9Wcu0Q28XGTnX0MWlzUIg8g
WVbc1k7Rpv1fLWnmH0fiycB28/GWHZ6eVmEDxDwdOH2sVDT8IPyS00VWq5Sd7PJW8uqPrlsDaepr
QpWxiXk6XwAjbBdQw8I0fBz/+pdz9ecrxw77q5IMgiSZf37wtAe+GHhXl7ymV6OzOBMscFXi+0DH
P1pxHrxBkHH5VO9RiTJb8MVkiieVy9EmnApaFgcyRRxpzCmXdteMezrvNuHUeHeVlWq7YWjqr8wT
QZlnRQ6Vw5YZTu6JfEXZFZVZKPQJ7yWDXekRwa2tKPbNEnJorBdOdVAtq6JgnOlg8viNLmStWVJh
w4sYIPGzkPRzu2i4LNerI/QcOg2hDk7IcB3nVrKSRQdPcSLsAQivEeBlntlN3ZxJ1g1kgtVdFaph
JZa56KbNh4iYRPq+dZbQMyEfCa6nbuso//zwB2GNF3gDCdaMy7+tjHquUkAqjtIvsOAFJysDAETR
TtqawiQ697MmWlmRPqESuRZkN+7CbwlaMoGfA63Va8fdUlxIZqWAkTNT5zoJruMJXncirZB1E5vK
7MUH0kIBmcj/v80mxq8oDypv9PcKrsQd6vWAsseLzDmfu4UjFDzBdCouAgzt5va7Bk0ejL9pSzF0
eOurDMTE7EO0lKUlYP0J923qh5m3U097yGc27pgv0WQb0nUvA1Y9Bhr1Q4PH5Qn36PoSTHcNBpBz
qONTqQVYtoa434/SYQDQhZ+mVkpq4f7GhdSH4FhD1p+u8zUv006e2isjBBwy1TOHONnx9DAxaErj
eXaQB5f8S9Bh6EZL5PcgmnckkzBkycDsUAQmgz1qRE2ijioGeEpFWfCP2OYfXUeZvxKbH8mWBz10
v3WmyBz1vQwsvB6dzrxPZCUeVX/MZ71ljPxy6faCzHRzKseuf9Ajf+hUHgZbCJ/FOgqtXWsUz+QA
BAPS7JzuZzYdWRS+M8uKd+zJ0vKw//fUa2AzEWqmF3GlxL9FlYkIWVhMeuVBXJAEyWnfmlwaIqzX
/0yz8dIw2MAWeIVg+oge1Lp03nSGyRQRq2pt013MccuULpoQM2CLiVaPfB8OEiuN+tWfvqxs+cIS
kSDW9BFNOuuaooJi3FVrgpeZjN8r4VOsxU9cg93ksa0jkwhKwb4OJAcN0pQylbBtlH5V5I9zU40G
stXlESwV8saVDeoyivSvaO72FuD0DdlVQt+jyko/dp5fymmUfbJVIhKmbqVZXI2/0eXFcL8orjgU
9C1XimjCoumS74ogAc6+3zXSkahieWVLoYX3tQpe/GrVzlABYZXGKRhld2xr/bSjDnSTxNyKjDcU
zUh0toaTCbexxAB3ZaVLwOTQlTptDrD0cDw1+UUdwYXwfmkrKhJKRDi/zVVczM5iApAzjlfQL/gx
UlYGh1F2ckcsCb+UofIwcn+qJgdVagWh7gkwN5Ev2HcvHaf4Elwxt8k2isPvKl1uvYvznVCw1y7F
AXzIElOiAd//NrNpfnEXmLOWALEWZUMy+92H8gyUDs/c3QivUakY+Rq9EU4BilS9CNz8T6iv4hHD
poet8I1qOFMVtG8GzSAqCW/POJXT/0FQa+i3nGAf8/HGpqALIlv282cXOF+zvuOlhh3YGOw0n7Y8
CSPFo3rN1awDlEe9tBjTZzqC5WjsqdXq4aUXBSqPJ1k5QEnZYjqeWTI9bzQjVNl67GW33ScYU1qM
fAjtBySvztuW7XYUmSePMDnqDNb0xLTH9cwfT/EE+qp9PObIZYLtBcnZBthWpNa3y54W53xL74bj
l5fd7JW1Y5monTmOxDJhJikxHgWwVVifUw5MppMiS+W2WlTjAW5g/xSE9Om4nqIegNdvfJ+s12t2
yoxvrEfVMpdC+HoW8Ze6E/sd3P8d5Wo1ef4gvCyKOX61P9R9rZg7+5pQVP4lp2QZR9xTnVPeiGUc
07Y0MZj71a2C5CC2wLlnEFg2biGfvhqNvwfYnzrTS/LFZeyxTcfPnPMV8Ylxvw2Nqp6QFzGXOK7B
E+WiO/Sq9dCZ+hWg/FNdQqnyjJErtyIniuXIJ+/NhxzMteNkYXYJIcElwBqluYW/dEepsnyS8wYN
F/unMKpVJDEm2dbSOllJ6pWoZktAtOnUm/anctVsf8FUqI2GrU38Fb0nOvGeTlOuKPrRjPGuME7K
PlBxiS8ouoAYX3kgs6xvrGArAlIJfsvXlckA9IA0v4D3M2W1F2LgV3QssETBVjIVQxJPjzWOBr2B
QvKV1ltDFOgr79+8GBG4CPHQxJI5NHYTN7pLEj7gw1UnUBwoLpapLfOlIAXG9ImA7xINI7SozM4h
zhQRIJzIUTuFLm2MbykawYkh4Ht0765GVPOhULckSa7VuDiglHPMe5WEi3tFyQiAbCcK1G4xe448
z0ELnzxLtntoTL6YySr5ckQ9s6B/g9/0EssWCjOWT0bzJYdzWMLiMpUbcKWjrFgsEb0JuoQPe9ka
q6wzjsQz3neTGVq07bd4tMwc/ao4z/XEHZQDmmqeQa08QjVTE9GzudjgEsSg8BJAA+OkR2lJxG0f
XSmMuIsvK8OpYwTa9a4iwkKaIeCxcasP9tzpsfznThxDUKEIN45wp4v3HCYQu8rj+qP17bwGjW9V
bv0wHhpjEHsVx7FWE1QvMGijCq1EVQvNJyx8QJjXegn7wEBArD0X3l7SLLjwc/AOSTWo9oHhShIt
RovYGbikoscYoZMftYm82UxMN2JyXuXj4RWdpS5exEXu7TaKPqhUn441yppOkt5DRWgQ0L5LiXKI
aZ9DxNShyE3Wbphjc9txfXBpteTA4IT7OPnzoDBxPgkaC4HOOb4On4nCE4923ZBnbLza2eULjAYt
uHKlVB6TnU2VQktGbdTPKVAD1OltL+qm3HcrmOgilYH/rQZ7FootAXJj4lLKUxHYfiwZmS7e3ASV
qdMhH843Nmw2Va5YgZIO/3iR2ipv9pBiBWEm0i24dyoF2ve8p7gzSIiSHAWjdoWL3DG1kCBEIZcy
7xjCAi05j3D9TUdRqQTFr03Tn+GFVkSybVheNqtQEknazx1xWOqDszeSsIZS1U3LgpOIJk5zGDSw
qaln3A7T2xxBEI2Tc3YTf/RNN5ug+XTTNV2ECy/mX4U2g9Ea54dAoGutQ5HJL6OU7zIOCUYYEwFv
vDdV4RyIRRnaEdelC8vPWuksLeoDh6Z3zgP/AdUu5mrFO/q7kelKbOk1fFcl6gQzGN2bCYNGHo2r
89MYAXi+MP7RU1NzR5DpVFwMLlRodNysgeiM7WjO2yLy1Vv15FU8CsZ56P3E7vePmPsjFwbUQz1r
b+qx+vyN1Ahth1T/KygQFrxD1iCv5aWIR95X/oN47CfWPN6TYT2FOS2/shlrU9rp2xjuLffxZSHz
P1OmPYmKqva4wgtntk5G+DNRxWu95oUXafL/d1mnUhHC2GDFAcaCT0p8SDRBGy8TOUGuqx6FwWL2
9IFhHHECevqfJYheRBNHLfEZtn4062LgG9qIcPzQdaabE1Xaid/rP7GbnA6fM/vXmiOj9AvRmJEy
3aWVRnvyRwHD+FSZJj+eX1T2fxRt6vRlN7zFCvn6lMgUfV/vN8rqWF7wOGFOyjTLb63c8aPL64tE
mOL6r1KmAkmFnfndbwGYGE11bWCGw0mZ6nHdY4vVKr7HY5A3amhg1QO+tcdLfiMfZ15vNoS7CfBI
APXBK3NwZx2oxV37FhJ9ui1GrZHy4Dj2KN50v5Mc2t9TynvtVipGfYq9xKdHo4u7wuFHaiQ2h0GQ
Ff+qGXANXCrPefDCp1AR5HnSjvWxiR2H3Dek7Ag7njtbLqoYe+4hfiPOFoTelJr4jDjV2B6MpGEy
BQbSMQXHImuVSF+r1EKGLvt17EQ112wAKgDSaR+jDznovKhoh3JR4k1DRvTw/LFT+5r4ftTdD+t+
Tkv2E0N8M7I/nD+xV5KsxGZtcQso8oiA8ic6cM2e7SHXvQ7twO+wErOS+BIFa9dKbfNFGq48HZZT
ABZbA96lrraJiNap1hZErclxVuXV2KxOKJek/506onQ9/0eUnqgrw4wjtdZ+z0/hO43Vns5xxmwA
H/yeOSDyCvbDkDZ/vzBYIKzhb1RIehvAeYtTTm02jfOc9x9t/f1YkSzHXLdF/q3F8iQ696NdUUp+
SQ7xgMDpZTJh2J9x0nz7SgcR72awBqu9CISgAAl/RgRxXwy5T8AhT5nG2ms/qYOK2mZHqDbuckxu
CXnXpyj73PmZpnTu3NfYGP9z06D8wZGlBLjmfxrtXb/nq6kE28AiLP1DJaWlMLs5o7gm2jbY4GfE
wgBZ3EB8FePJkArarjoImUfNZAQ8WJDOlVPG5k+gq2NgRdXWd46toBckAcJdSidw1ZOQxSQ5n2V7
HVo2gkXRRI4xrIdx3ADIwG4bVENKUeSjx49oLZWrOHAjQWFjy15Jxn/pns0YWHzLBMmJmc6K/1Tk
VTirMZG7xw4ce4ck2+aPhSVPTpKNkdRoibsd/hNXysAf+Ym46D6wEs4g1+RgBNKMKzwsWVT8YLe9
tqhR15rJWxylxNOhRiv8b1BgTkFWsVydjrW+J9l6u119oLxxWCl1G9ygSoboDZhcqGrxaL/qOUyi
m2VeuMAvUkA4A7M3bmww5NgN5aCVuM2tEs/m1c2CptzKIEemdtqyPwBixnJ4Ps50xiXFqSM+eLmv
rUPDxNluYHV9GoOIc9qNblxTvMuvjMlt2dhBwUDa+wHT+3iZ2+mmnxrUmOMXmuwaZ/u3d3uvnPwQ
yW5yjTQN5f74Ueq2AQKskZenz4D7ff4O0epIwiNxQ1XTDCIsezHsQ0xqF7CB2NaIB5bWXJixd/Ri
0UsC07Pd3lTTMM2xXjtmPdEWg+qVIzNe0v2VGaVwI38kAv5I7ucHc0QFuYI050kAuovgFTWPo7Sh
P1zEW429FsnrFK/7qrAhJ4DBjccXkhaYuyTP3z5BN9q+9P9YtcaYd28j3WKnRaj5zOY/U/43ho85
fz3uZoYwRZ4Jso5Ct7U6KnzKmztulsAcgWDHg/5t7S0gEpR0McIv/i5btlDlL1IaCYVvYOJMDhtX
pRBLca6HitDTVlhjfzjHSlKCSa3rd/hcXH3xKOGKIUCa/7vCS5ayuaw0ivEl+Rv7UWAjfTgQ00RM
RRWEainljb6rzBSxAIlBxhn8TCEAqZeNm7lCoRrQyS44qvU85/M/vWheOpKsDGLMceFI5cvvv3EP
KyUt/L58TEHktlnX1iIU3mzRL73raT4DY5UlWAUpwmBTz/7a1cwMz4I/Mlj2kP2+KqYKHHK5vkFd
JeghmHHROFe3H08nndjky7HZmPZcWz7SsLBX4v3wb5bP2dXFOB5zmUAYY9uv+nZBvqmHuWe7Dcgv
L6o5Qizl0MAHaqE5Iy0y5BQB3NsCF8195+ZcZvYXz/sOoHwwF8aJGvkX99Z92vUljDB1tJoQkp2H
tVS19InXVFNUQHHLgl9O9+L8lPTzkGUqBkU1523CEZoc0pa+ahorf255luRyj8SLKhFE8hLgGawz
0X0EVa5IylgV/ARYvRcElVPmsDv2mR7QJBHjagCwHMlF480Hp9PEhWU4ppiKlHpbSOJoQ8wt+7P9
BerblapteS5fflmaBao6I4Xgl70UVJyFeLLRqsE8C7/GGF1TUs3QhWvUfUWMKpePub4ehfkoXEs/
sbPeMhhO9I2Ygc9lVKOu9mTloLECOF6DGP6CLJNuaftnVjCFsfb83XimksZUc/mL2kWTJsKkhonL
2yLcuWqa08imxjaTSti4tscYwYVsJ63sBM6bPZv1wdOMnKBEsXM+XstnH/ZZj8dBl+tskAigq8Hq
DNLpr+zKVDh7uq+RipP3iez9gejxowKjQ9LwWyPrqj9TLZjFEKKJktvf4kj6e6EHxO2aIiH6JfHd
AUev65UM+u9XSH0CeGmbtuUswxsMaHk1tTUP3/Le5/WP27HbplsygKqNLo/1lP5gg44W8nE8Rjt/
lDxkbJas2wj0vtov64z6ULKEJYeY+qA70cBuOz2CIumE3qCYo5z1j99Lntord9p94QNRy1FL5laI
KHh4f6WlBC1HGDtMVh6FU6hlWWNTog4qg/IfMq+kDmkxlxVCjWZmUz/592VMWzAAoAFMuvO452sD
8tV4I96CDQAYe6FeYS7OOIxO8YdSc/v6ZQfAPkU6oOVd83+ubHxOl1Q1BqL3Qm7hiuLf6kU0ojTb
2hkBuZHUWQxSIyBghrU0T0lyyUHurJDo6L2eO6PEXvaT/jFaLUZ61sOG+gz4emb90NiTD3XNsAxV
NEVm80ChYHP7+cozigYAaSmTeeMlOuLO2yxGPALjkiVcizAH7zc/hU3Y7FKv+29sBXKqOCkKNRnP
eZ4lvYgBPPP9+WJFQiJA0KNAo11M9llrDIAfQX1Hvbx6O7tP2KXlg+T2WVSGDIXkEHEo9UbBXyhU
KTcEjBYXDKMsuLAFCZWG0RAZU5+2OAB7sMhhwE/skcgzv8MmJZcNWotyt2LsAgOvbn58WWpa8JJ3
80I32EOd7LeHacC1BBvE9hevPYesiFvjK4xL1XBHSrlr4SCTNDwrHklebnuFdvKHlXFKKXhlN+x9
1QZieCHrzuJcifX8InO0/f8jCtMjme4IcLMAr/v/Yt7pn8jwlH9fVxt3U0LAMBYWd78lKt4dr/s5
OmTENEt8OEwGmCOQ7qOTaH+rszlmPKNiB0RSA5ckkD31KlCuKfA/5yM7QBVrZK7etyYuLNXRj/r7
iQCg94kjIDKGJ32O4ZmNvfPe+ThClyrDfCIhwM3zWVuNNSQtXC0oq11CWG9x10kT4AgrGCm7yEuX
Lcs+QyVgg0qiLD6zMFOhqs6GMXCclK0Q6Yl4teqLf9LSBmNrDxokJf0koNNy+lxUGqoz60CRhkOM
3Uj2N8nwSkADVoA7v4lLAjTPsU+F/tvf6uj0NkHaqULJNo5QVa9ppgxiV9Fd/hVGr7GTG8qEuNMY
rdw4gxTMbtIcWXEdcXLvKQgH7DZiQrdaoJHK59CckbmdAcJMcg8T4PrKDmPbZ0/uOmkBdnh9+8UT
OUHuMa0+EJVjdhSvU5yXytTiYqwfLz14+bUMnjEi/JuL6u49sErVCAL+DhL0rPOsEYSjzzdWas9N
6wIK6dTJ4W3bPCojmoP/CGxJmRx6aNZFYNVXuSajaPXZHv8ktaZEo++c4jUK5pTkr8Nm/3d2AGMg
lDwROU146+ChIDcZQKeD79PYrecKE6NglxRzg6NwvC0o2BhjGROwx9qtsK32/+KIiEUcfsOmNI6t
Y2rUUZxNWZB3bL6FHDWQAnf/qPTn0ZzbnAfI381IMRZLwvQo5pTDeETL6ehN9zB1EYFCS/IlXjfn
QD/kZ5iyA6qNBWIVU53BNNFgLvn55f4AaGejwsIAykDYRgQc6TgLVjWBCKKoaxiimoekSyqQTvPV
U2xQufYaeGDf5ZIY4duUWTjI/bYU6SGaIDf+SW/7gI0/5AAhKvbBOSpkzDyIhIIeXSCw/LgcUZgh
JFJ0OGhsur5E6pf1n+8obJQnSuZ5CXUfrtRUGQMlMd+KORrr5eyN2rnB+Pnn2jqlzbfqkf4XGgG9
x8CdVZa0hjjkeVPs9zuLLYeCczUKwpDvzxMPeNH0VPmRv4xQu6dofzI+OIDM65NzbWeSFMuH7nmt
MbXxokpd9hhStEqhAbXpzahweqldFIZdyeUzXrQ/Sf5xeUlL5E4dKbMKL3ahm2WbMdJKB3gnKe2e
yOuaelFr0aDAh9PtbrmLZHuG1r0TxYyxtb8hmALYAOqv5oX03GFW9fwapYPSeroe8E25QwsukBuA
De6511iiWOgoK0wuRwkTtMANJRbjLzjZRNu7+rziKzGmkenQgOru3BSQvDjKfn6b8Iq5BNqOlqpo
Y2A+PKwg4HFM77y5LrTXBJPaeuWEh8EUNHTcTB6T2FdWM0TRkFD2quCWv7DLcvOB4c9sWpHoadgV
XeAEmCue6/mxu2xHDquDVGqd5B8b+hbo600QVxU0d6sdKAIAxrxEiUxjPwNlFBz+OA4deTE5OiEM
y6UWstOHgGETbdreIUR1RQC4nrm+5Z9TQwif5a5r5Zen/d/m3Wz6HMKr5hPgWZihfm3kr80J6KUB
VIvsnmWJAjtBSUR5/u9dGyo7zcKQu7u5gjwNv2YGyb6MMZWc1GEsjl/D8oTAsqMd5JjePp1uH24z
8fDbfe58Vx04Hgy3cQEifI4OVsLn03eie04zQet1uhrlQJzJ9f0Gjfu7bfhiCpIeLUsAcZnoq9W/
J01oHED67iE3P+t14T2iq6emt7DiZMW6horCSWx3LmEDpcn/ff28Azk0loNORgl5JKAR8A1ogRcF
LUavo5rU+qux9z0NC1NdkweL7iLPFh9qiD/yKDFMY8sUotikemQe61CmJ2nQk0MZHrngu4zyUcdf
9Y+x9J/pa/AKn1sKE3gCiLQMpvNJbE1X5wDy11tDiqE94ibl/OTDcxdJUvXvPOgexDgChnvcvSOd
+qePo88ftE/SYDjg1StYJaUzML14xE0Kc5FzXAfiHdN2dDFyy24JROWjzJuRp7mh5Vs2TawnC6ai
X8mGpthPV0zd2wRKaWKajOEnEpPGiQaruKZwu+Mg0iKgq/fNq3w8X6hqqvCYwpoLf5517A1hyVJw
cg1fLpgfctrTmeXJ2MBDOiIoY/f3/oGxs8N10h8jXP7hT6wnwGI061Ui4L3ml7lMQE9SEjBuRmFp
hgo9FjT2ux+GpnKzRmNYkzv5BYe6QLMPqAIJ2e+EraPy9mmGTzTxIJolngOJXOOqDJBAfAcRCPXY
SyP2yisjiMf3XKC8DEgkIphzSKC8+sMqHB2D8XXPOAL9qxwdqnxhc0JpKJLQRKxfPQPfVViitb1/
MRvDzkHPkgEumDlKhkXBzXAU8ebWnXOE3j/Vjne5NK7+jE/BEBxcMdgMbrZ6MOkn9GVPplpQiNE2
piB9wDhxQzdSZE1jU+Lxz1cZO/WoMnN6begJWMeCAS2Ur7DGwu6Rur3IG3I7/mHlx8xxxqCP8A6k
2hSa9/5jvQhrwY/Jde+DF5rcnasZ9r1RsWQmxt6ggKK5mOIbI1Cb6iOtrNPIFATYnydujW4UsZMU
UULcGFIF4VuSPW8HEXwP5wra+Ptb/EhOii9exjQiWCqs1v7CTvT7k+rB7ByoKpe20V5NrI3HYESL
W8XgRA/mDxsQw7HbZ4ocan4WMYkI9f5SLt+tDU7VEVCMyd/SmBx3FWIQP2pyVfGZBl/RGTz5SeD6
JtwBa5OxBbrHZ8XOSGAiaSJUWwWyLzlkxuToRxqGy/HR/gDlCjFJuW2WbefkDk2+e4mrrpSBMeru
iz1Sakmqn7MRXkKsA63McZFzUNaSFE6dDejXpuUPLiTVTsZxs5L0YmmvmhSPpf14Krg/KLEuP8dI
vcdK/Brh14MXfHxXOBHvyPDcBQlfiT3JUqRVhf1hI7zfXyuZJATIp70mUQijMuPGbWgU0OXQxVNQ
Jo+r4KcGQMuvWVN6k9Y8fq4PdaAq94ijsh4oMzhozhPvkI0yXN1yEeHq1VauWtFM5qjKg+kJnNQ1
Xt4+sPDkaj021gBNRxXEZOIwa/DHb8R6i90NTPaIGx3vTEjXnfRO9aIpFwpogIPhEKJshIC94kmB
Zfu5MIo1VV/vmDvxCnQH5prxW5sGwhi5WIzXvYYvYCCiCZt4pgrC85chofHVkhMSwTbkWi7rimcU
/DBKWJcnWYwJqUytc4+02qh2tuKIWQsngPGdTw7eaan9Zzlfk8v2No/0kFb6ay2famfpg3AvM9Mk
rp+Ad6Zam7tu5mTgvoSwSH4SSj5txFQ+tAm44WJbkcBA615+W/ND88CbSaRN1r6f2wyqAj6ZUj0d
hrQNwrLE6DRRlUI9YHKBxqBsgS2nb1SyObBvPAAyjW3/T7oWmTAa3IQnzeG28EIERcP3Zkutbj1L
Nb7maO6BMegCbWTSoyPDBt3VhKz1uOQdEUA4Bjt1tuxYWqbEe8Vw6oHasAe6y8KYxW7mlJmegu0p
q5tbdAGvBgFyPo2GUyNtaHRZtsNa8rWXDg/vF6r74p277e3Yta/UAQRAPkj7EBjzKpaWMggegomf
4Dl7nMslE8CaFO2yaN3SbbNST1utdKIC0zjnb5wrLgHy/NgbfyCnE+HqadN8+0XFAAXmqb2Lj/bU
Buq4pwd9CM9COS8zeLamYwdd3xESgExwyqIDY2GNVUTx8IOL496zGTkUpoal2ZA82lb6vOyfdBbj
diua6NhlbLGIfnOC92mzSN3JIpMcbc2Mw01ATeQ1S99C5tlz2Lh/CJvocORO3PKM5MzY3ZE9rpr3
C5unxTKrpy9WFdOr5knip3uiPLSWDOjUaMpMfc4ti/c7hR0tBWVgIFntDS8RzzkvwZnPB+fedy8s
9qgRRTaVgpTX/qNwDZRAXwj6KlNdOd2OrXX0UVajxsZf1bOMT4J8iaBMzBTxWMN5rt1nVvpoktfE
freJoFJ+EB2gh49ZvZJRYJ1vk7epdzSNbrZUD7C90UA3R7kWJvMZ59s4FIweYFfLhKM5zvXhXOxC
irplO1epYJYk2TPHchOd7P6+z1hjwBvalNM7dwcgjBQnkY/kQcxGsYMgV2iQ305QwErY3i8l8AYx
rlcWp5z5v6XMD8eYQBfV+u4begY0cEbDVWI+Ogzhksh+v4EPzsXIG4MU91gPaD6PLMkwyiNIyvHN
AmJ7u5q8Vx9fd2z63juZxIpw5AIxu+g8LK8B75kPp98LslK04UwI1aSxqoG4t00LNFUExSsyatkf
0JRMc9V/P11ZIH2qn03/Z0q5KesudwbzxglzGH29p+jMSOg2xMM2xrBx693blVtaVKDmiGHUXIif
Cq0ihUH1/aP7VKC5+re48NbCRO6F974iijWHKfPljvoFDh9ICQTUMUTouGlzyOq+uK6xm4IfAKdz
wJCWhDd+06RXldPtcoA+Zk9vQWXKByw2vRvVFbxW6Ki9cw8Aikzj++OsrT4gr0iLqZsgYomG8Fdz
aBfDFbxiC2RLkKpgE3MsTwlMCtDhcJVRCBwYPgLf3CoUPwMWPU+9KHlxOqTPL6GnyLWsOB/7vklK
yvwjAlgK1DkCmy8ZeXE9AhBHJOmGxRq1gi9XIatzO9bCxLrrjX0yapBNJSvfyIVTqrmo6oZyvAsi
omxgyuAw5QfDJ6GlVhsi/ZgJjNnHPl7pbAMhlFHV/c7tainMcteOnLIfDfqfTvDBjMd4MdnOLzaE
cdBtqBj2HDPMSCiPoo9379kWDOddAKqJl5b9Il50owgRzk+GomDBLB+WpqqYQwYLUPN2aELi8+aY
SLLphR+uZvIEvPru0eEPs6c5sGpKfV5yjZAGJw9XyrrqNR8/qpFSPuvBbegOdHgWEAcVsoDvhCLa
dQzOsCSYtxGWEXl1D71v8EkFuJsupW+2Rdr9f4aUcsZnjaqUDhS0HlESNGvmrQoZf1P95D8lNu3c
iEl3caiQNI7N/sKb4mcqZGOyAVmplf4c97wbWkWtM5hfEykNd1Zz+LZ583F8z7MsPT7ujUykonu9
fTlQkN/ix0nIppwk563xPkSpt+umQKyrleXoVieFetRCm8FWOagi4x85/QDna5JAb4THlA7mhCwl
1CiQS8V6Twtfstxc7PygNI85Xm+QJUu7cYleJqWAnyGPweC7XIB/BxpiCPiJsYuMjS58jD3jT6g+
t9IqncH3pdy3mfLu+l9HjG7j3IB0wIB5OK4K9MKHmr8EPatrQK+9+pQaldlDZ40f8l1g1tYU6goG
B9YQaV7eIW0ky1gGDmRIGO05dH9t6wadHLL3pC2+aMm+xVsaEMNZ5XI4S0dojwtRyA9wIN8wqKCC
UoTD+xtiURI/pxcgrEgK4a9VIKjDRe3NylcUZ2Io10WotUzhlYFWxGWj+ZVJnUsbLD0jQkGay1U3
rrLDcC5qB+KfaxTYXYaNghbs8/TmMovCbbaB4Jh6yAj5dz/9GeCB80opsKuIq965pECAM0mhyzD3
WLaojGqHKBMmk4JANUPPzLAq14NpamImqe4pgdt41fmeCs1PfBJiUwB5mXjAGKa4vuMnQ82t2bSe
XGzzBwuxZg66Mvri0TYbg8tio1dOoWIgoS1TBaaagT1z8imHBZZGxpuANayZjHpoDkTDbbW6g5JP
BNDrZs5IAfFdXW8AetC9zcnBmm4OZnrHyZvvFFTsMEKW6vSEXVRUqyI0huPGJsgkf1wmJQsKOmXu
whJ21tIsiUeniwjxHxoNCJVKO9zRODrn4pPmwwom/3AEsHPejvkVFVqyE2I3cT+GFZzdPbPqF5pg
xulUvOa973Xg8h3BVts/8bWHasvRdUVxENLXS1HqgvLHnoJSOyuNcN2C5eYLNCXAUxVFQpvAu6Yb
b+jWfn5jQLxx1ZP0BqjddKp0N+oxBepN3W3fERiJpC2/Q5iUP86KLWRlRADp5SPj0dioVOusrpLe
gG3QtfbogdycWmLFXuam4mJ2d+QZvJ791VRSBxGwH6/1Lmd9yd6Wq+3d1ahnNwdrB8a/tVpCw927
JiajCTPywxazjiIc93n2MqeioBHSB1Chi3XW2FYB2TRwMlaedTHN4cP5qu83treG1Fd22xcqkdh2
eM1pAKPAgA9OxcPnsX+po2pI83iHSzIVaV6qYxyt0oe22UEgUvjitAKTwmnD+0etT3w4UKAUE3Sn
W4tFOUUc1ntmAeqt6auXF9s/PlAbKQPoB4D/Ef13nKM+OZ5IQZSV0qb2/ZcmibnB2X1uGaTMHpQM
CcXWe+z72FpVjZ3rC0yju7h7+7g2Hc8jKocLATqmQPkNHj4eIwprllgSBP3b8OEBV+mWg7m1TkyO
tTXmNF0BoXHu3+s2dUpFiAZLyVwAfuZW7QMF22J7SNThTy++f5rC6sUCqC8ZCsabVqeD+Akj1olX
L2jXzb32wSAJVC1Sgd9NbCebM65KvibsekZOP/z4sK30vAywYAiUCmtAp3Otjku0XVouo4ur1TTD
dHBR5NnObRT5eETBK4u8AiFqRI++QJkw5Y2KsJjCU9/ZNYWyYnzdJ53hx6ZIxJMpL9PzCYFrb5fz
DZBlm1i7XkSVX4zUWM+CeJBCYu3xI41fmaFEQYAxq66uEHQ+WH2u8WzOP1th4gG1WItbKNb/EtcZ
P7Wt8isSg7JBcY5uUM+v8NRQFGRnCfFdZPhgTB8IsxN/uTDtzcOaB6mN5plchMqaq6FtUROVelN3
bssGKui49QvkqQ7IeDx59PzneANplYiPPxWA1c4vSc+vAl986ABMFdyB3ByB2fCZtbyNjwzLFJr6
ll07TornKcLy3LOsYD9AKZJsLdxgYqRsjJnuN6WzQeROCtKIowzmHEk1nj1uuPu02mW0usjN9BjL
InH9KWPBwNo8NsLB2sp3S64Qg9HVs3yr6cnMuKqzEgiXR/5P3ZmnOJ0ob/Thim20bLtbeITYIwJB
1xr4BbGDrTrvVq+jG/ZsI9pL0cRqtZINP0EZBk/lJsuTSbCZnX1LmSOsIPNBaxYvHkDJ8vQ7I9G1
cIWCnnrQ3N0652dCxXd0VKpYXkVC3cnDuIXphYZOmjrRQqqPhhDdyfHqyFztIqAu+yzelnkOVuyc
04m4wDCKpgtvM0cQguRhefq87Bbwka9V+5pEk8rlvHmviz/bNwQxxHK7zVoCACnLfXp/IB1dH0Vm
15Mn2UUN54PKLMJ4bMvBzlWpMM85w3TUcrgv8vLL8NE88K6o2/z50UvKyXIHC6gLM2d1hiytqazT
5xyM9je+07Kmale6bs0EXngOtRpst3JQrAEmKpCjN0JF5lkqd+4EEW+WEXdhv0M5evg4f8Ftwr+K
iGpzcMfUNql2cavzOWj41SQuxkZUYvxsswEH/kUFp6XK9bMR7Ihl2GhmcocM9KRpwedL3M5gXU7H
s+/6sTFopta2co5LKwYdMbZblRT6G8iEsikwOLhWWi/AGrin/s9DIVlQqCLWj2jXJqzx5KSd58i6
/sJmGBliEjtiv88nnnry1hb8X9qItWQtfM3NM05aBQRF61IB9QEuY+fhUGkrG8kgoiToGYhJ7Ep8
nu79cPIQ0i4GT1JrmaTWOniHitEamZQFfx7sO4ev+N3BNtnGtSVRUbSjKRzvbS13qZqOVZZ1Sb73
BaKkiRMum3zSZq3TVegPXyMcMB9o6GN/Xdt3zJ8RpdIgu9T8iOW1aBjmUFWJqY75E+/c/KL0b07p
EQj7nnfu1pli7QMF2xM5F9vO3k54Mjvl56zHJ7QD9slB5p8B7P3FkntmMTRoWHsu9z6/OruMn8IQ
Ay4NcH2iFNdwfMFQ/3ZmlMsjp5K6JFxVc49g+3S57whQ9NWiHF3FD6PsobNKSYS103L/ZQNoCAkA
x3EBjkhlqko49vks8nRYiRQK5yBpEiEDuOONEV6nVT2R8ZWQReJPLfjLdhxGnZHsqNmV6BR1Z3jx
St7RAocy9ppNLPxJ5RMBnH03LCVVuh/6j8zDdhGHxmSm+LQffsnkihS/Lnc47LTDaca/xEYmyKED
3w1/btvy4sP5DtxKfLHE6mdPf+9li2c5WpLSld72PVjMb6W4rSycBliDBCLa1/M+DLCtAqu0YQQA
gI9QNK1UcWu7qaeiRtllVo/WdIqwEhvyMwWL+kVWWAv+hJZf3z3qUKZcw9QSNZvmtsByc/AMNSeP
dT5Gvd77tVQj9BcZlC7rxDzh6mKNzX4Emv5DaRhTmKA0Mz0a1gN6L/HsGYM69iF6nq3bDK443X+B
Ad6f9FT+9D0/+9ym2XktY7L3WIXqis9UjUX8EY4LbROQ0uyOUtG5WuTnryr4l8NESEgv5kjoDHe7
5Qp9H0td5Ge+zanxOo+duNmx2ePQVwJUso9dwLG0Eaia/XODbyF+FPOc9WApqLfqzbz3KTI7S4z4
xSt/3bu9KrMNUglXmbbsx6jNOO+1koKQIc57FuAB3Wk6ZDDXOHpY0LbqOmadGxgoZrOcaZWHsqbH
x/J3Z+Zu2i8eHXlwRlilTn6NNmz0PATjjs43wV6N6HxLGW69aEhnjFO6Wl1xyh9MaOiDn/3H5Xmt
V0iFcpwZCmSbN7lkJObdlzwrXGZrJcFBsrXymQqzBtNjhhrIRbswwR1UvOiyKBE2BL31/TyTIeIw
9Ul6Li7UBanMiZHtjY4+66fmG96BAydfGDku7+liAMaJ8hCLKZNLkS44CSJiHm6CwoqDmbPfn6iF
IPGpqq+ma1WWOZz8zdcLUeWUE65adH85x2Dr51djNs7r6cVHZoAy9Xfvz/znw/ojdWtPyOyDLAQY
ouukKqgnZ9gex/c4zTWe1VQT8SLbfkaOTKwXCVhvv+Pq9vCMN9fShIDjVoDdjnI63OnnTjksX3sP
NBeazA6AFpsug7hnwrL+5SofdK+4+sk+Zv7qRUgHuI2blHLM1Q8HPP/reg7Wew5dvh4f31fYViHx
886mOsMqVRgZeuFPE+hA0gKKfljmrekY86J1gvXFyq6y1aTguYpgf5Ebxtkp/pj/hBoBBFMjbhNZ
ffNx+ibO5NjjJiLZvX1jUUJMuC8Wfc5wr+cBvKbx+8txokHgQPzbGeavI0poe7Tp0q+ehWq9N3eF
DQYgXucqL69gNtHO0CYoFC5e0ZrTBZTy3RG4Th0XT/JqxxwehxJT3+H4zb6BW7fGkHfEtkALjIFv
ODmgefCfGmOQEczTIxeF4cfSo8TTsCrjIRj50R4/xdWdjl1YXsMRBjZNsHJc9ao/Y9KLZeDAyTnC
qJZrsvBgW7GMp11lIBc5t4HkmOJ5V38sfPL3+aNUqgYlp3vYcJkaLQ4sg0DsDnbnTCir9kCx+SK4
71gKWTCKJGmqKdIHnrzhC9ZmKBmZfYLG+ewpPx9VnddxhTfZsqxn9Ng4LzGJf2Bz41FZz4VFvP3z
3axrjCUnmpO+lE7xX8QnlR4z7yITi4mLojWFmkvIM3YtqJgT0Ahcz8rqkte0u3K3zGDy26+8UQex
6R09Hgt9Xs5AEfQ6shST9oF2bbUCIhVr1gvWYvl6rbvoFgJA9WqdqtBFSFBEpIW0U0x83s4bKUII
qT/89iKl2Ub+qnM4oLSkJHla5tKbxPmcFRVYBlANAExsP7LYxgIQFMAZbkVdD1d4bz7YcBxHbN4r
HdVsWeH4wjQTmJu8Z2TnxAGQXfcTgLeDnE5gx8ynOwO/5pdA8f1L2FLJ+o8/eN+84pD1QQVXfRE0
uhAl2ijnataF7eFDQhls4FxlfaXySEJ0JCTcoLIBapFF+yBEnBw70lB4SbueE/4uyr15qS5SgydJ
3FUEdhC18aO2/gb5kd9Ue3gRhdBHVIp4mkBPLbyiyXhUcMbllaMKfYPyBGtAptEyCMpDir3Ck0FU
aHdVVj5c0o5TmeDWkek+Rt/JanlDfvBAWewLlPac6o3ITMGTmrT+4uHHsAlsSyX3jsGdfhI3K6RY
ysEBaCkNesstT4v4kBnXGK5jqjmQdIp7GrUDLnPiG1oZYgEAu6NQfhItCFpbAGjXisU3T2h8jmr1
BTCrHCpLKOYo8zigJQrxOBweZWb57yBL3ZfBYgdWuaxoFfygfM05+MP7RoFkOFegVXwKQHB2Y4VA
jpOBiIkjtTjCv6igdNRfgA+uyjH6Tzay8yirgh6rW2ctbtcj/rkhyzyHjEtj7OAE8xmS47ChsSL8
wiBYWHTdLzKFp9sHU1Ya4eZrvUl+nDZDOEFwRf7fzWRww4Rc0lvik6xYYYyFU0R4uuCWXYIcD9Wz
FBiXenSJ9UqUema/rlZrkYMavAb+mdv53g7Ss2P1X8sSxF917kHqjqGcHARTgK255e3zs4mMfjAa
nSvIz+Z/0WgQ4K39h37ph48omEzh/D0RFxkEhW4SUDpl9jBKXlB7XFrrBawb6MAmghABO+SOfJjl
8yPbqaLioG/8IPVGS4PW8ku4xUiCU9MrP8fUUBFQDCu3smM4KDCqgi3qXoCDwAS+K+ovCEgvCoCB
99x7/xlePmWEh89xD7Zer5gRr9dxTbdzl0AkjbcMzYhG9emWRjxVk029ip4SzCLJMKFy+0sJkuH2
SJmJWAEnvxOFd7Dv7giMiv4VQmZqPrB6DoPnMxpesFB/4ZVwpwQRfjflJFtuLFIe7n+m1WPmdORk
+1HqSJpKzLeh8P/8SAxCZ1BAyLWFHMT7FekXwtEwyuKd7ZgqbF2VkZXcj+6rP+OQLby8zEXt3VYB
GMg29E8DngDpjsKFB1KMYqW/iS5oI1Ssl9Z4JSeS8A7lqPsAIbuxfWsAvbrN7gJfSKFyc+bykV+w
QR50kT+fB9SwzHqWBEkybwdUz820+tX84efDf7mu6AoOYN0zjikjDTlV9iz60BP6Am1GJbUw1V5q
E+mqMH8BsNnY6pBwdDJF2qoDIbelJ5W0x6CEzQBbunB+E6AZZaPnwybPPByHKSU3yzCq+/kMtsGi
iK2VcnOqxGtKL/xJ+wCFQWEt2em/jaz2hIeav3V0FsmU5b1lQiyQdiZnvGXoI4gADqulgEW65U6g
ZUpB4Adb4cdY7Pe2fntavyqPb5bjRJiW8qORAVSEYKDgMl0vz+0GY9XEWsu0Y4TOqm/DFmpSqlam
8RN41vTwlmLb3ZKyXoZ5IJGl+T0bK25YRxYVpvqkvloIafvG3uYxLyvzUPLtLCS+MAj8e4GcFCU3
AcnYrI9Iqrj0tLk4kzyuWaqyC2gfSGc324x898Dv+mBS8TM7bf3WaTBb+bfNZ8PK+xP6IxoI5hNG
32fu6ILsk0VEf0Jt1rXuJeDWgSZi8yd4xYxi6mynSPy/urvbGse/QMzeRjuOEfo8g5LWQyuZsAP+
aR5RlxGwBVtLKHqUq4X6AKSdn/5iY+tfD2stUGLDNY+6XRN3FNfXUfzbSXcF8dcC25ypCyh/sb28
E4dOoFA+f0Er4qP43n4kuJ097J2jlKWzLyp/sVSQwPZ8MOTQENp23zOEqwIHh/VWSrXC/bl8F0Cr
M/7GjKqcvU30veFxlJQFLye+jC+1FN6OOSnOx1NwgjRWm8TQ1q6nUU75RW7fxnjwJ6JoBuYfS+qr
8YhRBAhpIbHBagrttsAGsTcBzmlhAE1KUJzqSMQMdAACXil/jHWH8LrTuRUMX6cCQLqi52CfgmN6
Ak5ANpILJ6wtcl0OJybaad9q5YKTb8XTYegSEqFqCWpOn1kHaaon7HhEteclUXkuCicfIzmfoaGH
XgQ4fcrzeLFncA+zI4W820D6kT3bwUFZ/zdRSwy2+/e4GPmPka10CHfrkCI17CnZ779lJlaD/3dt
xOeDaL/C/n31dSkslao+n6gP/jYOhEgHCuJmQEhMQRLtayk/bVRakH3aJp1YHPgp3evSNpak7k3M
14vCPnPnaZN19C5udBLpqDMpeHjTqBUIQSLD3gVUCNJWY+eEzCziXwCEL/kQ19fIM+Yzc33aqw20
DxwXc41cx5S5ZCRUA/yEr/7jP9I1ytCLXoE4wwB38Mu5eMM6KKHJdGL0EO1rZaPwU8sELSPB+J7B
EeELgSDO4FkXTWaumSL+rGYWWOzEgf0nMgFvTMtaTg0GPtfDf+MPmbGi6kqsifSOnxKbaxMHPsiK
oZr7qBd4DEa1aQu62ypZNOUoWJjIlS2wCEK4gKM2b86o1gaaL0RIuVXjrOhmjgxTRgnii1GCrXjl
B/xQnYA8Png1sMEkFRTAIkuLR0+kTIEtwYGR8BwLqJMRq1n+JaFm+S/yXlWvU+wsEkT75cJ/Cvet
GQgRAwr4gQXDDSc6iD7x1Wyj5mlrm6gKOK6k1rJQdfI+qc1mjQIL278LVrNeWf/F+x1hMUBw9XGw
TqJMiXv9ArbBmtAmIr30Cbc8HVSuwOzMRCgu0zOv68Uhx7WULGQpNqJNlpdxAxTwODnIxOJ+9Tn4
UPvD1cnkwy3sBZnewgsECQeFmshWXK+ykaXYWWVk7VGczhPZp3yKQQFDo1eLMHP0u/2U7xfWaJmF
OX1nP6LKtPWPpoSUzurADb0UXoRLCSKqIAvbpFDMaUCY7y6cZrlGSnlLg43rQyoYZX/BYkHX5N1/
nnZHvUqZj00ABVI3jYvx08BG9CqQeRP9G5zqpxzpe9rxqTLtfNlmDUVDsshQJJpITKiz80q7SBXR
4uXQtiBQ5Kii61QBQQEZvPI0cGKOyFimgm8KL2LzlyR8biCcGcRf3YnSKlev4vVpO/sEYEGyPV0W
4or3nCWQpjqkqPTRf3XQaYxC+AxRTz9Bw1yG5v6pDd6jDi5vUUn6i7UUHVKLZMITC3068JePQyjC
tllH150FaFys8DeclcK1HPU4xs1sheLw46R7uKO8cvpPMcDAHZIW3e8Ad/OOt9vAhF15PtnUKIhQ
xONW6DqebmhqVp7P2PJQnRCaZlO93Fg8uC2QqWIPpFJvlRXQCHFioPS5Q2e7VOektOWEvqZwiQcQ
LouXbEet6N2Bjb9/8dx3lNkfyP8NrMyFaFNge6TpjPt7uF/kt4Sp7EzTcjc5JT+64QUR1C9mGmFs
MBjlgrNS4MwH6c1u77oJ8Ac6tKdqYftCG3e6+5fDf8xediatpFFwTOfZsjHDJ3B1whXYVRbwBg19
KlVSFi5oj9AcCESYYSbMpNgmMN8X2l9NoI/Bhkh96sZLAVo482dw+UvAAQ2FQcO7QY8TNr4Xg9Zw
IlvVqsQPqpVddno5/ScDGrNYlJOijfiZ7MLWP6iiNMogHQb3KHCkhj2//XHqDzDKNoTImdIzSZF9
usf+NEzIh24kvROmV3LZygvWx9CSy1FE8aoaGDLq4WQrtW3LBy85bXLaNDHh5Tu0zFoYbcIegFxy
XPT8FU4NTlN3TgEySo71ZKiMg+teZqJQrux0wkdATyi0TZtsbLACcndbKK7FbJg5I44pAiK8/ADl
Ni5dgiBZyeXdP8t3/vY/aW2QLqLsDF8Bt2pEYF8LOFxd1VSXMkZ7UWgGvS8wFLlBpuc+5+hLMW+/
fQV48Siok2K6f9JRboO0ZRldOOh9/CsUNyfYxTB5py2Sg/xUgR+ICFJOuqcIYnI4o21T7BxuhTob
8X2ADjJBg50PmyiTznuemNh2EcuBkK/QNfMhWHflxJEEnS8bpKa6cnLpyFCM3SPcj2pme2sDA2bq
GYoId+Cpe7FK15mjWmLbgryI0VcYOSIOeZUAIsy01XKQTkX+onHsLN62drHVpw3q+cpYi0bMLUAY
GqaKo/gmxbk/i6aAeg89x1vMx54sLZFJ72zaSh6EXpCG4exXCsR8he2YLdAtcy+ESuXCFfsHDr0U
3D5k8iNQUlBWGVVAFHKYfGvYvDh+jZLqrH3dm22OO7gBHx7RNFsszI2DWzADQJ2y+ArMqaR6+El6
25FQS/6dyP9dBDMSuCxXCLoE1PS8MX7Njz7odmckr6MI7UuWLQld/Flori8+1cBAG+pXJNaVuv9+
dFj/gWRXsrzKq2iQs65obpoIiP+VRMU/ZsU+aSqQRsiy02IDqt0j7PO1qZpdEj9Akrt1336juqlg
T2C0WHtLJ2ue1aIXsgWAtogDpcaFel5CJbaTUnLwJyP07VB+Fr44/SZAwJuDG+ScjnsSj3i41m+d
C37/f6jrklKLrkUDv2z6maTeRnhbz0Ea1luBKog7ZN/6IxLN4A2CTIWy1tFtsNVBPs+e3kK9TJRl
T7ABuPKl3cL81hKYcx5Lx4rkPUH+4pDFSPfXoA7H43wNT6p1R4mVY+GqQo4/LGXdbk5yjgGNNL69
0p4TH+KYxXFf+wYO37lJCyCm2NPftGPoyaLwqTeS6ennCAb5LzJWCEP4+rUC7t7TZjeWXjbKjZnS
b0lHVhU35SxctA6PoB4r8GbWGRIskF2mCleO0kb9p4LrbSVS9SqTNWH0Zz0LXzJQ0vAsgHwN9u/F
+Y+i4I9RJdRaDC82cgLnGAIS3VBC0SdBbNtq4BIayUonZVtWABd+2B5AHfjkubBpVfTOhySkUjAJ
89Z7G6tLHxG898FNBqDQGEXWUxoNBgnId63Yu3Mn5n1mZv94xB2moSnb/Ya0CagM+NkhwePG8lR4
gnuiRq8pVOOUJJOzOCOjDTFuSs0Swwy0TkE/GLPhV439uzgATIwNLjrd5IMnrbb2IIyt0JN3fj5a
ExHWfYuah3068+88xnCs9LAfFHbKLPJZxvSOzSe6hONqNQsyU8qqmfN2gX5pj7WkK/Y6npB9OZD0
wo1PZDQ5YJPopFK9V/2YmTJxNOSjr+fSdSZd3qKZaLB8OejIouztqpY/6U0RSe/7t6itA7/i1DzP
S4JQHN6DRKfAH+omCVgua1B8cCOBnWsVOb+ZDnKKIvMdfayAJBKPI64C0/gpVYXY4Tvu3wCVjV03
qqqJnl7cK/x7EpDevY8yd6QlTjJtpP9UalyKcsAiymXyDcGuGrJAO0lKYnBpHyzb8cCMcCdtGZDU
R6iEPryc5ItDsXrg+K4ZOIpQtmr6qucTBvSNm1f042OptzP2/ouj/LzVqv+HgmVs5K0iAIDrcN6N
gxCvy2uT/WwGqF/4YFwH0S+lnNcDuoILt2ONtDPWgxoCbxyqwcD5D2dlSL7snUpk1p+Hg0/Yd8E/
Uu5JmQZWWLMqS1MH2sAAzbPb+wmDieYj9O8flxfiouWDzPhbSWRjOgou5KbgPPqCaHToJGYwsaNy
bg6fUfaOkhb6wAehM21OcKZcK1WgHJp1yEYUHPZ64AzT3H4fW8aXcDM2xshYlnxjS2ZQmnY9cNCj
BFJbYsVGu2ROzjNc6feZa312iMNmI4oV3b6IqJ3YDNpMq1zIFHynk7togxgzPCvHAMf/HRajGX/7
bJ76PHgVrmb8Z4fd4eKagChdRcBSTQjhYgaj+eoNopFfysH8IduaNsoj/Py2LzzvL2xH6WHPK8Jk
nUzdUICkPQWUYcsMPAl0T8h6PUOf070BP9EWOZlSWfa9BFu25bW5xtcLrtcrzM9TIacYy2i7UCZU
nS9VZ3kbI1D/+nLXGHNSRseq+U6VyfBEvmLM0DwicWHVDvcXcqu0HIBSpJ8HotRhNykNtK/9ZCix
yvjeB2Ci4lfHCmBUw5YSThbFYsudIs0PydrbB39+BGynbu67vEGAb61QbDY0et1A0W+PtC6Gaf3G
HlnYVER6mpHw1inrwClBFunINuJwIzhIRvBokwXAeiVsoFdRrqj4pP2kin9Tic60dwDhkZ9ZYFij
Y09Cz5YrGg67909fYrY6OQNkpofXm3bzKGv7upaKqiz8CvcSXignuV/WVIf3/CRdn8Ok4XIpAVZx
yLA9vCB5mYYlP5F3VDhigVJsL8R6g81Uoba8BU+WIQdv5IgyGIzS9HASrvfvRe19Ls6lR3Cs93QV
C0cWhtyDRiZ+kt63jpdxetjDbfUMojXhWcnfN2x+Va1CGHD2P7+UUB6vRqmi13CCnRAXZjoZdDST
XG0BDZGcfeYwEm19qntnLsstX584JvXHkS/yPYDhikd9fdNEZOrqBe+F5/LWYniLNnsEHRQ1X2OO
tA+cjmCYAU19LO+a+8BLsxAQHfUpcY/gpnyVfb2o0oyPe5LYGLpuaxG6on4ejkp7YyKKgCpJjWAe
BuP01LZYAmLrkVYds6oT++fW3Kvwj4Yp3Z2ftdiEXKJ59n+5ltbSj9HNIIeYBy5ktsi0vgN2zNUR
DFp9zzcyj56DpKI6t07D0XRmxxn95+9BR2ImTW09VfYFuYLAXyKx0ojdQyNa0pG8S5rZx2mUTkYv
lyK0DVUfhIUs1I5pZ7hIkX07iEKYNzJfMQK2J+kXsW1GOFkkhKueMpE+0NkPmvVULrRyv0MfaMml
0XsjZPdOrRXMeOQ99d21pCwOWUhcFqlKWNfLARKkfa5/jeW1ovdxL7SLTBnCS6/gR2F9EQvSerKG
z3WUzOroE/6IKy1G6LD+KxIT+VRrRjdytdBhPSVnIBAWLGUY122hJ8K8m+tNiofvquHgve4vrVjb
QssUQTtuqvxuJ9GtBexwbQi6VeVSHvwNfTiXbD6Xc3T3ht5i0CqUtO2z+C8nKQeUiW7kUfv/cEZ+
hfdF1COuUfI+87yrqcRyqkb+JZsMFMQY4t8h1RUdCGhLaBlHk9QLXtTEKRavqQ/3TtjfpX/UnZuc
1UpOvK0tKcLOrTGex3kd+BrFM9+4UmjXGRXQBZTaJjeni9tWKztIucYCQ87ycVhtfurqE64Ip3UV
pUXjxPCl3IeqWSwUnifQR7xWCovdB2+RaGPm9++rtKOFVWKSC1HVbq6NZnji7IiPONBMxdA8pJbR
s4oBxVft/OZqF2KOyX6Ldz/Gl8rXgjjfldChyES/PW7IX9WRZQGsGKeSbEAs7pHdCHlpjeOgSueO
IBL7qeldk6yBY8JVgpS3R8JO0Rb8Llz+oVg27M3o/GGTxljQZuZI5LZ5QKvHGUITF39CuUfB9AOy
IoWsoVl56qwFLMjk59ouGCFwjg6dWX1iLY1AoSDTC/bHarBnr0M6GGfyu5KfDjRoDi7Rw1Eq443L
dvJnXJYTWrNPBZA+H+12oV/SbFlyDDMeiyeM9+hgcHCFv4THKLyRf3nx5KE2sRRgQtNeUTbRKKoL
lAY7LZjkNNKThTYOboGD6iTby9zvbHfFSUX+SHRZaS2EMYvjHYigEDODV/KHpNx5/ZIrmVqIiQ1C
1Zx9jT5luPAIf+32swytFouNr+p/RN2tKSVxcD1n9F/VXU58nJa6uOz0JXops/Upy+O1ypC0oOer
xZaJhpCqeEvR9J83CCMhzOEL4XVgX949y7szveFaRfZ9i62SBEGNmpZLR4ED1LZsc+qUHwVIPbvW
lC74Z97OmhrxiZSIQ93htsZO1fY90iJ6tvY/kjcZa0x22v7KJimFD3PY7xDjyS6rDZBIsbPhgsyj
P8SHXhnpm7qyYy/9TFeYZnc+7rbDU5FBEcK7Udx8Cv/SKSvMrLTeDzZAsG0jljxdfci5v8gKt8q6
JT7sB7WOUqrUAHVzd/KEhntwoIcMIJmD1g9kKeQZBY6x8nHb7nNKeFgvhe+YSsfaeLMIJThQ03+x
eJjU3RuQ2+F4myBwNf+UXESHCnl8NvqsBozm8UdymG5G5ta8rNMlz0OlhdINTFmgB3JWu1bi0A6p
jvgG6M0vsxdeFrlD4cOj7QgjcBM4ZA+ahR/uoYJ/VUkAXeINgWeXWrAjfKVDqNUxrMwP1A9G3r/q
31OItdWzS4f96rZYxSR9k8Wz2JEnbri45DjSUJKANCvzvvH6wXIkSNfbuPlFHQgRD5AAUWvSpfXn
QTH5xKqVh3D9270RQ/ozKba5DhBBEJTRNJitB+7JCdHDrst6ZnnQ9SDH/cj12QaGACv9uwJ8WAn8
hHFLvY2XrQu/8b/W1UHjCBTDNcWS8crrhApDuK6Dpv66jIgetN5Bwee0HLZKYdvs7vV6zkUwdc8x
t6EOITTAlnu0Y2LqmAYnWZb1UXHT0hKA1u3kxQudz+FQyg7kt4dL656INc011yjTU5xABe5XhGkU
a4qiWzUNbmEKNwj5DeJNE1/YNPEfPBQ8rUWV2263Rst86nKagei3QRcHIe1ZoqEDE5pcFCnccxOz
3+xwVoZ6ngCXXrjYPxH7AZCpiwd2rxkUAnM2pW/Qrx+nX3uTBJ61DEm+rFY+ZpzaIuYwgmqZOGjn
2m4nwHJ8REc+uBNWIZHIu97uzxGd9usL1kR5tqZEqzQJUCK9uyYBPQJMJPL86sgcNVCOZou6r3KI
pUqAl4CqMeQ4yH4CHtj8Wg3mxoohiMlbMvZezNQZ/G8CLg3eQQ6jQLdr+kFSMXNYySUDS/FiNW2o
5GIV0mCe9gEyvoHaJW/GPpyXoqtxQiO0KvHaPYYi3sSMo/S1QaCyWuwWkDEjdexoXpO+cEKAU8bU
Jeh1YRS5J93hOokcNZ38jCeMWr1u6CDhGaYk0hU9g4W2CFbuG+3ZkrS1h34DzhHSd1mf5mZ3zYay
eMy5qM4hclch0Xg2xdICQrCEUWiCmYJ8NCpKf5YNMktM7/AZdQbC7EJ2MvoV5rKW7ch8PzOBr5DE
GzfLq7N1gzf7bp929AQpLsdFV+x0iwX7f0kHQ/0mpJ5UQ/j9dPerXZvWv/1PQHe04m8cEILzV+9P
oTCkMXi2K1JNfMs+ZJYNgxpODzBU9Ks+ZfrqTBe2fSbzsv6O/3WUMQdmvImQLU4SNQbv4hqAjmEr
C8YcARppeG2Q2BCRiKsW3cFiQXNEci7aIz9mGKILu0Qumf7qD/LX59vFpNkfU1yn7HxmiFK27sNH
baFsZ2DG85fPBVIdcxDHe1waeAjM1O7nogLmB8hT1sSn3mEB5or2t+nJtIJU2GRGVO7st9GtjJtW
rOO5VG2k5rFB+TTE7a0lLGyRCS3PIF8wOV0yJSVJE5lGj8yahDLdWjvoI1Q6IT+ndaxbCDGE3HT9
rVBoxZSL7MASW3miiM7VhDZlPo8D0kdSLFbF+lYfkice5vg7odvKuKb2P3PazsIIgZeeOwHIhsTu
NBejL0qrnwsxdMXDADd/pdB0djjXEbG7AwGpWCspWTYcrLvaU9bdXhTlXEyAursOuUqWEO86LBEW
/y0z0E+RE5QIe/6YjnHX2u6lFrEsZ9J15Ebq4si6tpF6mYMEn2cycM9oTHu7e+c62QIcm2pwDeeg
eX89AnAfb/8VVgRWOdr2AqWW0iZ9ec+fORfChdW3OIJoRtT/gMAlbb/TR/pPsVgJxOSvfHL/baum
cKZx4i8jwq9efS8Onm5Iad9eiTNOr0ohW/042zZeY8mRhgwdds9YT9drV2jQVvYo48maQEBQjwvw
VKWdj7VD3mvNSSormGVeHSedVa32wQcWb2j4u8GEaaNhRQOnc6av22a2tk3TLtT3gC0gWcPvSlrc
xcnQdpTjPsWxCKWB8PlUxXbq31xiA/Mn/LsNtIzF8dilq5Aks0Z45WrAXN84wlvPyscRYQoSt1Yf
wJYIEbdFozktXNtF0yi8GDlZ49uvqolV3WP/lEMVxUKuRC8Qdd3YfNRXWODGJwi+jZlfgc4aLdoD
YRaPdcTMrgVh6M3Kox4V8Ptu13mMVNh+Inz2wadovtMyFbMS8hbx+oqWWmInefSLtvqu67EjWvvt
KJpCMt1bjmbe3NzJZ8T7wtJ0O5S4JBRgZYiqzJZymTcJEwv3XSCDl81+OnKo2ZPgvQ0PAIAZLCKM
RAipRCxr0y4upfyQaFhLq0w6Q4Iyx94OeQNUSbJAUYciTIR0UVp4JAga3htHCo7bdTkUvb0eTgnW
nlUz0UCxbXNvTi5l+IHLFr4OCtP+Vav2sq9jUkd7xTIBQ8MUiZTEfyP0kTGsJtZh21W4wpfGaTvI
DxBfxUanvCn2YzX/IVUe68bHaSth4c6qqMOhQVwJseCkMQkZcXh+qSVR59Gnrz+oMQQpgr6CHZxQ
wFY2xfPx545vgRLx3uPZM7Ff36IjBjIurUqHyIsNr+n6GkkjVL+fG3hFf8ldGS/89oSOxt5cEQEb
t5JMBQJ/2VzHN5GlD70lTSg/eNetqyQUlA0sUt+J8gwx+Vz3hh2ngTDJ9RHa8egUm4vc0QB8E7ha
sdjIUbqpwScFwB9281nczpeSzlPGMsMkORU2QcfPeuWu92skQE/yUjc7qZVO4oADu20k3RMzvSjx
RzlsjNKt6H9yBiHjZv56BVfkNWAZJo8+79Vw83uu6WCJJggerbfswrWGi+YnaJWQ5aXg7kc+O69G
q7IFuJkI+5wGmPP1JkaiyDLIIxSU62dRX1gz6Y6oL2fPBFJdWBxrpIQeSBAvmqFWv5MjUiekqLd1
ZfLXAy8hYVC7nQOlpXg0jwnjcumCGPjC+Ce12lWsV7tmhIL41DWztx5FhG+0yh0g4NSobVMbVur/
oorCKEduELOZdZzsvmW+5CmIqU0CdlLATOoCtsGQBbmtqCZ/9nQSDYTfPrQFAT15BTsxLlEXzb3E
DbMG4zVcMajD26Dubu6m5lYAjBP8F5c8wqwgYa2xY2dOP+tVEKXmUzj8fdQENnzOF7ruSTT2J0zt
E0LDg0ehwUMhAgU9yPGcCeBcTNxdSwH+uJNgVHJPcNI8kuRrhC1S2smBVzhzwOmy1tRRxrpAMBGZ
PHgRxQXoRuD1jZjCEGE3xo2jd8BXRLDk+wWjb0gXY2P33FutsF7F5eVahFGlLmTzcKzTTYuOgXU+
OQKNAm3ijQhr8Yfv5uJHDpnxyURchtGExKku3/L8emfA6clC1cJT/XnlYwvGLXyRKxGJaXU+wy0Z
V2e47HybTbEO8hsFFSzbwkX55QK+wu0YVxXEF0A2n4Zec3eEQz8D00uDGRPzxjVo0dwapNqqfo89
y/s7LNIVPtT8JWg2lpWEqzGR/CDo5/AR5poLR1edg/aHKX8+94O6bvv71lrv6u03HydwBPJ/2wAo
WAEjdxQ713w3281MmWkSrvnzRzBz2vBDPpoSAyW81VuJN+bi3fWW8tYt+HetIBWAsCSag/3o89Rl
3SrmspF3TtYVb303yf3uZGy7N3xP0mXpeOEwElZ2n5aeqSRSXdTcUiBL2K0u07KVztB5rgxGKFm0
0pXhI5yDlAa9NH6RiQ==
`protect end_protected
