-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HVKQNle6ZkpMjsCLqpG6zom0rf6uAbivbzBWT/8oVBiw9nPt9iPmwpcqYvYKZNtqxBh6+AvNnqZO
WaoN4c0Gbhx8kSRvKeyDQhhZX2hO0nGVgApTT9wQqjmPHfCLNzSIhrLtpNEfRYOLOmzS56sjhSXc
U6SsbOaeQ9zeZP1+1adv6WwiMgCYpwCLh9RnCitW7U2BzOQ/M7ZJ7HX6triXNOEo30STAkV+mKO5
XmxRUU+a/A0yKpMyy/IOeHUzSaXVAn+LEoQCgGz8L0Q8ql/VaOKmhQFadNHf+IOA0akChrTyleT3
U9rUXcCCr4vMAW7H29pklCn3jvlK9wfIpEdkHQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4832)
`protect data_block
48R9L7IUq7Mxcdc8S3AJcYnGftk2QZkxbJAuDs40gtBLqg5tDqSbj3Gsq0a4hP4EZ3ji5AOCkikP
o/v8NJLhGrwevOvQYIXGzVCy+EbQ9tR9/Oq9MKqs8KixKPok4rSHe148WGCWUL1OLXqE85gGDAYR
Yu/bzsjMwetzB1vhDtwI67+ujveVoAwY4wzbypLFgUarDQABa63kYHp9NpcBGl/nQQcGBagha1F2
9cKOBNmBOj3axDDiAt6X6pUuxkyvUZibBMjsKSIAHxDXVzBeB5G/qpkq88/0xcJ4r8NcXKJDU5qF
kD/VvlEytbNlQKdBSDBXWu09OKq1Ega/HVjcJMe4JwFxyJv31BO6glkWsSytuXOvlkpdPyCGrdN6
jrEVb1UzqRcjmuroVlmdGllOZ/42Q0kns5XoS6q34/+pPuyppMVxRLBk/87yVfttCPFYBy8oQ76N
AG57fHFQEhgm+4VPVv8QdrjUbac1me/o1MJKiV5jKIlzM32IYkHnIr+6SfPltOCXeU+aVjXBA1RA
d0jK7TydLfqeuml0RJDcoho5YFSJOqEo+u2a9wUXwklWXByk5nIwvqHxgEDfjT8FGaqsJDU7g2e6
cr+Vismp6SKWlsNccuwvjOyRxbx3pBVUtRq2zDlY+yx0nTIlzviEMr0hSADjfIAHKrx0o5iGuMyZ
NoFuYH86jfYY3kA2GasJXKSOTnnIfdKQc/l4D88WkoM+TBdziHzZ/5KiwTI11T2HzCos6cgK3GmX
eAYaVTZZNfbeQDEJxXSsRaUmUAdYJmiRlZSiZ79y4lqIeWsBC/pZMviTq9IyMa0OTUqCbjusyUiQ
8fL2LQeeZwur2pHmp+DPmr9kuJOsDNWIYJBTfUgnt32fx5a3m8OmZkJdD92WAn/Qv5G4YcImu2Hx
pJuVHjhobu0AqUJMzNR5wvw6bSiwZ8pWFmTC3oAL7TZzl0wC/XlMMg9rbZH1i5Otl2oxnepTaKeX
x7lD6eIvfIocftWfCvhQKroyel1VWpEj4kA6bOowwaEqDRULHA1d7orTmKZESc9tFDyo2LpxYIZK
rd/8f3N+/MRRKJpXBBDswgA5gqoc5/Xx81iw6HQElgZDkDHBMCbCOxxldbB3/8nUshakJt30XfAL
LQ6cFARaeqA7VRRQj8ypUhSQmVlp9xXzqTR8i2/39KIrC5yW7ZeNGOldMsi9HRJ740fPsSn8sQ3B
8OpeB+qyND6+lg6KmtBgFaEjk4XNf2FaupPMQQm//Y/b/NQjju1G4vbG6Glw6YCb2/wO4cjnBJoB
oO1wYkHE1KVRhoGrE4HsjXFiu/kTf5W5RRpgzOM+o2uuyUjtnl3lmrCNArk9DWTXEBqVzZkvGhNw
LbWnWQV4bKxJdwEQ/zUt5B9mhGvCoN8fmlTbUbxwayjAIBHO2HufxJIf0ak42hno54oc4WS9fgZR
kLsZZI1HH3WCvP53LUXy2yNVJ3OfRqYvSjrkuTcglSBqSC17bjm4hQnCUNoJOAE3cjrVJCX9EM9V
9503wP+gV9Ahf4Uk1RnEWS+YjTTKJ2CWKRBOBsCqPKvH2zyzNSklAtJAlwwomZXtaW5R8AC6k30Y
CVyo4BFb2Cawt//672dk5twQVbvRd5+CTFs/hoLj0SE08sH9X8NEfq9/TMVYJ9J45/98/owdnbIm
JV4EjfjciDPcSZrZtqrloM49Vou5q8talFz/z4PpJzfL0p1IzLQBoumCY5hm3Fxh/GIJoJGsZVzn
XFiVZ/uz6UNe/nPYKKj9t0mloZ7/JL8yFIwQWIkwkeLIowWgCUI0aGlLzPdkmoom5e+vABhJ/jSx
7pI3p7Ri0nTDThwGbb9p96UIKIr1NfmZ5nhF+6N0Ki5B7oJrkzc3c+f7kAC6gBCK+yWArOQxcOA0
v8nmGQb/4z9ka6KnBJzscY64eDGDtd/NXyXRjo7UrJApLbCGAmr1vKMetV29rgi5uIv6H/Z2+VI7
hZ/Lv2pAeIxQwiBP8SwzV6S3o0CN8N3X39x2rYukL+MgOiPlAcGNYgluRIacR0oMehWgJ/IzyqxV
L1ZoPUO0dOmg4zwNL8/4xAbotWH36cAVbRfDkqfWYKJADGW+iIBYuKEx6A3QXZ4bOe2EqE5qPhrJ
LrNToDEnvhyHKvqKXI3RItTI+tAVcFtAyxJLJ+yaIMh+cWYEwQ+06oRaBa7md3nX/7VwMaERe+0M
jPDdL7WHSA1Jw+g52SnECKTIAwquqYUZlT7ZdDJBsTqIlWZk/099IRN0L02MBBhd2cUObjKOMXY6
3B6AvW1vbn2p++SvMnYc64PpnS0TkBoSS7bs86v/i7X9utf+75M8Z3xi0JbAN9L3pLaE9FMCAa9X
Ny5QrxIaHAxMnwyhTDbtvHSPXDtpnQj+sx3x4MvX8j/oFmnFaTt8Eqi3KIjB0LKeOYprS5Uk+Rt5
rFmNYToKH01Qp35Qsw7eQKbpuGrmUSjqdZM9xZSIoDEgZmQmXYLy+S5zWnp5YmjYp+YW1KEKk6d8
a8GV1pOSgtwcjitSJJfdfAOwT8Xp3AJAlywOSrxfJ679GSuuLje8cM19h8ajZEitOhN9p7O5B+k1
mueUa6V37JBHf4yt0JyaRsKo34Vj4cvR8oc0pYAhOEMTvzf+DKqnn/NHQ3DSLzp92zhFjvKH64x3
uf65XpM/EBkXdgYvd2Z/F6so7MdK89sZ2VCPQvdEJ53KKM3Kdw+8AXLRY1t4UUiK/CZzYP21da8Z
fCQVUZ46pIpoTc3+DrA39LGDL4miIicdc8/vrbZeHlT7fR7z4GUc8Gquf4VkMjewVUR+2F2Spscv
0rtrcFExxWDIfGFDjvJMYFjOuKmFcUBxu7xYlopTmOa+Su5y0ECdQwuUoQgKMaYKTfFw8TJDBmgi
M09JQbZGZ7M8f7F6sXAHJfr93Bd/FD3472UCunKrxMkqR7lVIOPnj18K5DpV6U6S04e8Kuqvzs/r
S6nzXK75AjbcyF4MDVFtyaNMy3l59LJ4LRdbFWAwlKJRTWrRd3h569Icu7LmYjaw+dugz9GvL+xd
2NSZTey38i0RB+CjWCOiVZQj3USEBrJq5UDScYWNqjf6C3ZO76KGYI+0mGJ88g7UaofxV/1pzHrE
X+Po+EWu7W3E+/h2M2qPSqY5nVIGUAsfG+HOK0VeRyeVMsipcx+uEWNhlmSgcGHr7KCcBZif4B2n
COQzaKqm44YZxuSpeguAMQriOAQ9jFooZnToZZJkd4ILRMklArv0blfIwAYqbPYi74vESy9dANJK
oB0nh/MB9+ybm3G3JcavqWX0gDzZk+kfneCWL/o21NUBhhvyfPkc5G/r7H+8UmGA8yL0TNtXD8LV
ocWfAiZOiKBChWR/gq8gaKlE/xOA0xR7QQPZRTYeZgHxPwBiDvkG24LsGnpiq4WZWElIyJ8D0eBL
qYTD4pzp0Ej8tbB4fS3r/7+rTFJXvLtr9sjAoIKqWA3Nv5rvb7ICdnDBrUcMYHCNBIC3HoCN/Rq0
rUOkCwtTqlEaImVBLn8c8EruZVGbpS8NUY19KyGdHEDvw3brPQxVpdo8nERsyQsvQnoQZIdvtM8q
0B9rxUDxVM2vIV1jltCy5TPPGe6NCczucUbNPYGt/jOAgHF7amu654IWuzvFf7ZFBpq3de1XooGs
2Ovw2Fmjmg+JPB/YtUCUe68A6pg5EAO6PWNyd7FQ9yy6VjQLI7IWzhALPF2IgP+ORXDGBIHW/q5M
MhR4H2E/jrC/8gK6BTjHadKj6yfjoEhqQYX02JY/wJJkCV+Qhkdx0Xtrgq9wd5+ojgB1ynMAc6Tb
73iPBU4QfSefEcFe3+/eRBL0KL5NYuk93DvT4YUsAj6cg5Vrw8cKdr7VT6NGEWYWl7lHN/Kz4jKN
bIDEkzEU6nrsukkVFFbt8B6JvBNsh/Cl7AhzBwqWHy+7p/ICQjpjoLZarSwREjn2Mn4VcQx7ZR5U
ANODB1/IRxqdWFdQc8kaYl2sEZjoEnwzftKvkFHX7yyW/ChxsFSv4/p8yHwj/bc0Jngfz0TSOpAL
u59Fz+dgksAE1LMC2xsVhRu/oCmbYAZ+WxIMnPwwJxk7awl1tUi2HAYkTKCPyzLWka9GPPLhUVZt
j+x7qs36r/FX7icORtF9LqCf9qzzDGShtzbh2qLkBocR2kCowUln96kgQm68Jo4amjxdYrVvHrjJ
ahkc8A6Ao3cVDGrKmvh9gSujsF1Ko828RhNmQM0juh+Vfw3okrBEeMy+0tSYZe/nm5UNG81X6tob
2aUpE5aFj+dcqY6fZsPdZXCeYC1065f9jIYnUh0XLQ6jS0nLVW+3uC99txk4Cc2x0FeT8pbsSehr
4TUv6mMAcI2QPOwTuEOkL4Y42f6u8uy3e29j/+7UxDCZPV+bQhq4kr5uLcjf8qiSnn/usWCLW2xx
/qPO14GqrPibx0IqxDrShcMA+c9OwCPcUI/xInVaj4TWm7kQmabQmJotyStdnEXWWyyRr/bZLhBv
QhnsD78JrpuVsuci7JX78Ps1drPzehLotdwO1gOao+nFqPTPTBpfIOtI6nN7G5AaEX1G/ZR1MZUP
hlaIU9Cm4XJ032j5p9AKWCueP7OkGIbqSY8wAl7h32zRIgBRS2spVr2g/QkUkHhxEa3RTSY4sSyu
1Prt0ocm+IPBFWRUynML/PbykIQDeadOsR/5G0tPwGND0lm2gi86iOK5mYkZHfaTPMmv6qf0FJ9m
Cr/Tq5hN/LsQMUQdwQsq+JUZCuGrEhFZ3wfz4QBJUt2LndrrAqIx7w9lBX6bq67K6V3eZE513PJ7
DqlwbQb9rwosqjpBK7Mn5SFVFP8Md1bIpVUo0s+RNtu1jXu2BEZsZufwfFN7Xp0LXpEw76h5c1Zo
iP2BnGIlPpgGcT/IOs6FZa/wFVwIGrCzC5hImnEtIdVdSIT1o9QruDaRGOIhieiNZSHJxFW/X+Bi
mQzuydqqSXC1jDuG9uoVx6kPLm4R0BSsecFp3ffSWE4vUWbXb2tlekAVv67fyK8+japg93paqPiC
9k1eIObVn61A2xj+/r7NJYVph1vXRs337Lg6WM3AIOEysPj3EP0IaR8gaungXLrT14ltt+wl/0NA
yAUrD6NvpgYUcjGZdbjuhNvA0I7Q9mlKlFrztt58XRsnfIXuTh3o88HEyDzF6o/cl5ztDqadDOMF
a+hHHha6+WQp/kJ0qwlGGuRkwGAi663iUZ8OfyFVIQOuuFkt1C4kW4EpDs8iO6rSMjj9T1txG91Q
QL8lTTWJrU/I1MReu+HOe1Mzi7mJmOXFqGgcg2LoGPQpGeIN3sqlMoZxHD8He6uerD7qNW3GjdGP
+n37w34l7awmAMqC0xCqG+l72+eWeewaVL+kz+bye47/pt1KKCFFzTajs2iMU6v01wKhiyjy9ilP
UEWV3YcfkiR0o3SUQRjt3NWLzL6v7GFWxbbskJZw8UBcgenwYGh9FDO1zekZvKS4i38AXCHrM7Ru
xiBA3ASPZhBim0VLoAsrGJnKFyFlB/ByiQd8VmLkC4GiGPQbJpC7aoLqx7AYOC6RW25F2U6SjQsT
jB2JE8wQcBE2bp+WhaPWK0SXvw+3RuS5RFTU9WSRf36fflxMffh4nm2UAafBhxST08JiOototAXm
DCwwQ4JMNrHExdl8N0eZW9VMr0uvOM7yBS55YbJ53pJSAEbwvZUyGudt04UTBRPRVfaEGsL/GAoE
GnLxYSyblQUs4nQqbMsW638ytRP+QZhK/Xa+wGz3UlXMC46T2z3hQeIgDiErZh+IbDYOSiJ1w/UZ
94CuenVawoB4MeRKThL5zcEycBHPgsVo0ukPIM/GXPm/BeTGj00bSjnUvbvhRAg4xD432OAQNhio
i6Q7UjDsfVCUgGjfB2Gajas8q/3/q2pAK24yPYn4lwojB9L54lgSkV70Kihl8SgizhN8wbEgUIAw
lsTtMlo0SobmqGluw81IokltfP++G6YowU8AfwztqZOK8zk+MjAkST3bW+3tMFY8bwZZjjOX/RNG
Ofe81FIiTJV8pXSdV3kCoTkOdzQwJZotv6IIUdy6dYsWKUkzi7MoIROLZFXck0bPDC7wpvbbkyHH
VWylDUn7KkkYwxvkjy4AycCJzX5nBi6wbTVqAfyw9fsmCfsjZx8xS8P/oCiSuMXcb9MgI8bT3aMS
9yiqI9KKMRoj5CMjUD8Fp+BfHj9JVkukAes2GWa1jguVUHygxs3uSLVTDAzhmbIz+ANiWEV+3sRh
TOZp7ghZJIp9oyhE6peeszVeCLJmh0bkCzoEdHzAxKecx0ZULAuhPFYBhDlgiVnB8McROnkoK8R8
1+eSETI6FFMAeEvfnBXhPQQX7el3XytPvWoYD2hMD4FfbF3NQzQJW+iWw15CJ3QyuEl0eWj4Ipzu
TYkLpokRM8+3gUnoRQLkM4qEBOOO8Gbm89xtl/XLqFIWM+M7tQz/Ctdvnm0=
`protect end_protected
