-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qEJ/8qf3P51kfXvBu8D57sRSRmeWwUfbw57dtJxPHUu1M0hhAlQlrPKmNJxcU18spwfk1o/BwA+P
o6vLJaHZelN7fsANM1MT8o4bfVRU6J14dBOzBLb2i4ovrP7P3W84/snRVXD50Qy5UCz7+p4syD4M
5rOR35RI9KWLZF+2N0MBK1XlHlsZ1o2d96H/L3fnYE30Q9k+OzQx7qqHufGXpBzs0RSspcUUikKL
t+sRQOdu1Byfw7MMlq8KvH+Pg9cH+YBYDtHM2JWxl9jzC+H7ZS96jjsC5VPYLxKGroA1P1fcQi85
RmzOtzk/7DqDpPj9djPSKIznXJfo+SZ8MBNWkQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8208)
`protect data_block
A54QDc6QRgxu7g9lRzpFndkdkkhKE9dFD0s3lcRi2VYl/uYfXd7Po+10YwNFwVCIe4S+zO9v+cQ4
NVl+Gmz76/FRApOkeq0XHUr/lQSnBBLJqF+BKeEzmztRti92ifTlI6++8Hm6LugWFZFk4h/tfkuY
StMzQ1H0N+IE9471epT/S8lJmI2jeP110+uxEjmajwmVguN1PdmNtlxyRrh6/4VySQd1Aa6GCLEe
Ux0m6/x0epT5S6v49vk+PBaqPGenhG3+0ViTirmtsaVWVKkHlzvTibjicfszb0d4jUfKBAOg8TWn
54zgUfFoVGeCfYplGxrQf8UtAvbapjbB4sNYUfnOy6fYxcW0LDM9uFMIxAJ+qpIiD4QA5FAEch/n
53D48kS2W92+TEj7jpPrUwjFnaB0Sqju9qWYu4PnLthY9bSzXNXGPimqmbZ7G1C9CSQeYZPMLt6o
i+yRSYL50JuJbVS/F7irciAWkdmXcXoNwgJiWZfqt/ChZYnH9b4CLwPo8Vfqzv96dY5ieKGZxPQm
os4SbFYIHmWE8IVRsNahtPJqwcq3PtOQfk0C2vA98aLkDUx9bHeeo9Jv10E5/51iqXFdNxDo0Wmc
FlSeiWM6dKoJSRk/+hsdUbGDPa0DDjxdiBo/Ge4wFkA+zyyErFfOXqReSQzjwapOPGnrx2wZGFhK
qddqSRCNFHrhU5SfSbwPMTdivQIb/gxf9bg11by4u9Jjoe3HB2ciqqnk8Givd9aWBjE4f4sZiJrD
t2tqLxvtqB/Uy0yKkvNLZXrDQ/xiIZ7wRdlepvqCpEx7ak02Ze7Tc17SjO3O9U7Kzx1QFEaFCJgP
dws6TzTdTTs8PFvcCqJ8UhpD+xLX1NaLPNXe/2H2pC1hYD44PmJ1AhySBAGZC/OD5isUk08cptmu
SBTovurYsWsuz7bKWMlnlQJPf4B2s8Z0bvBHr2PwA/Zprg92e6ZzTc/jjFMBPtGufZhuxN0yVNxe
u3zAzRTJfMDMT52pr4PgtYjG48D7V+C+EWFXvWBHLbYGpx2hvODbPvLgPAJdRTipTZa9Gc30TlJ0
NTAgM1q/RSfwZ8YKPduDY+VDna7Z+K+Pn9FlToxU9hKoC55B9o3kOjFF78MrO7jGPPykKrgaHPil
In+wmLaFXP50RNXK7gObLYO0PoQVaAQuAaxEfPh3rsH1hdzTSSTECCIMQJwX+ATaAViu7zii77VB
CHvaIqAU084VdWfolDD3QA2l8qbeDdkjzX84iYJDZfwFqGClQgEt2qwLOm8ctgFzVIbNQNm87XDw
8x1niRZe5BdFJHsuvOYf1Abkr/Ny81Kg41Nj0eGNN1Wqazhj6vP0rxovjxBLc0nBR7TkKnX3cPMB
2mYCdjP8LA17JZqokRpf5i+Pt8myQu/vigkApyVtGXRMibUbjCzi1keqWVSKtUjBkyhRjo8geVLg
0bivMPle6DRUUuKYOhlvyEJsAoUSSWt1mwK0KWEFmffcJsjVpQEoUfAr5o0jPbwb9BlFdSH7LJFs
G2vIa5Qlh1179HMplpF1Fnv9G3eI8x9tN4cIVgzGxfbYVNv2Y8PA817F6t6xJdoPjfVtjcg4ZTOF
SZqsfuLe5olk+qqPviEjvsAGH/bySQ6hQIy0UJUIH//gIcHGN6QeO35XLW22e0AwzKgxR4ifdYfL
3M1xO/YpwBUoqCcl6h/fVGBkMUlCC3Qyt3W2UFgstfWSDhHOBVLrpHRR6MSef5GZkTOjb++SWom2
b8q9M/OznKMWxNoAqKdgLXneKVf7/UN7PJ4DCvNDIlbp9eiIJMURAPOVOtMbZD90e+9iodww6WqM
Q/u82XpaP7/c1Ei3EP24o3vEQoafyzL6OYKPwJFvxKi4s+O675DTgakiBzS90VlxvK1uoFqGT5mn
kfAeQrHKOUQQHcH8ow7JFczZrB+XRm89ft386SFnb5/75hXXjkjLn8Sj33xJBlZ+mTy+YkAEm3zt
9tbd+rhlo7O0zGayXZKvBlOwVqe4ak+fVOPYDgVDWFs7vfT54Fou0MyxRwWXg7w5qmFujeA9Q6Ky
hplUB3ey/qry4kJezYB53JHUC+dp8U3lCF4d7tBTY8KBGsioaqUFKHfVNEh0XW8UNam87BGnzFRd
8ZIWqXVtcpvuiSEed4giOeXNLmLaleBAo1bJZRbNQvpucg64ZUPK+3Xs9Nimqm6FHbIpFJp5vcEC
t2nvBQk97YF7PWnzLt2hJXYIeaNsewn2R4hr6Xs3MqMekdgBgi4SPj1YLgeFfOAVy0yPRsJPGzPb
g8vYB8ZiEgudApWXP3ei6Dknd2bRl3DBZ9BMiQsQTx9DPTtVmO8DdvrvJEiwvO6VeD0gycyhMAbi
88nnVB9ZGnuuBkYi+K0LocBIJB7quNfZWpZXiEHjMMGepUg4hzQS8Q05ilSUJxIRWcK2THkTgX8d
B9J8dLACT8sSIXXwTLPAIEwzZCGPVSAfULwUnVKAfVyb/wz4V7IWmSAHGFNiUSi3C3RNbSXC567+
C+MoS05b9nOJe+SIJKnPflVUBO0aqOZedQ+5Z1P2phKbCZKs+ZIAkSj/Bo96YA7hERBQog8Qro8L
QxLyHCJ6BB1W7uKzhUKgK9RN4zyJAV87gjbQf1rGmRdnI+Y7OE8ZAmROBtVf1/6r0vRclIO7H/28
Q4PXPThtz2eCYzQKQuYYzISqz3qJVdJSF9PKxvK+FidTeBRFb68ouWO/x7eB4yrVkP+SeGxRV5W5
eBeGfWaKWZDSgEsUReQH5aEmD4Ji5EK0aCK80uM7TJHL5YWozgu3Qe3+zs+CXl0e4dF2OCFRbEWc
mWJXRHofnzFRBmxIpjed2AiGBCmYsSKxDSSURj6wBafOFDWfFntCaaucPGOAjL9OwO+WKjZdskpg
IbV/wsGf+UwzRUKKydvgFTS/ZSkxXqDTDVo6KNsBeCYIi5iYwL8vybyoYz+R0qIVX7f2/Lc4xRQE
LTru7j8Lq8GxSgFeY+oeEZQ0wa5P81+NdOxXg1H379kKXbSshppt856987HBM5T/Vj5BNpqjlWnY
u4H1ULkgmVerLk+SqrzQ5siqjspp/C+G8mzpqfmfKl6onun79KWvFayYu3M/3jwE7HhW17eo1QY4
VWUqNvTwz5aixMt9TXb6TnJMO8rzJhes/vT0AHtPJita08cSkEEhi8y0qENvnzet4plzMiJOAs/x
lE538gQ7KDRBIuTnQLUAVJJCGt7NhmvZvnvcH+Hu/xs9pb88M5e5qychB+5AWKaDIBeoJCYMqvIR
U+afWOz5umNsMp4pIpHQAQEMWhUPacwx7Me1XKMHyzhW9DjiNBizsE4GNZ1hFFrv+Q8k1CS+wMID
cp43gqTEW2qo2B+lGUs3QTZHutWveQxHpHs984rjQ+SFdLLosf8OLLMgSGRQEmqsDBVshfklvBkj
YPc/Eay1e9mzNk3EE3dwF8YSthBdQxnGCj8fy2h/9IAH3F6SpmWkDS+/k5CeJdahpRQ8stX0S+Ge
pCl2CKZAKkLfXK4nc2P1tg1jzQMWQFS3UFK23UjVN1sSg/4RsTaE2hPeGoU62dXP9Zs938hiQIAR
9thfwscr3yotCLRY85Bn62m3pEWfMUcYhK5aiBpLejXKga/7oiXx91jTvrFzFDLBDUyOEk8bpn5v
Goc4Nps9yUQS8LPrOmMJhUcCRgXhpbNFtCcva3qcowfy2YIk61RExVkN/VCyGhAt6xHBcRI1Jkbc
VXJP/oe9VdpVPzxALFiiHOWvSo2x46P45dzl/rFim+AzzLjVrv/+D4yYwNKOS5u4PdAW7VWSgVHI
odVgre7gY9EVGvmKYbb6Iwn+evI0m0hdp8ARRB/yDuTtAv2Zg4gGusXX7OCYI2AdUdkqoTqrNKiP
3eO+N+Xj04d+xzhCra/7foENsVPkZT3dgCt5603UZuMd/m/7QH+lJ0ldQmOUDspTrGSPszEWrFcu
TseEWJcgg8s02tbq7DVsJlOt6JPoUD0Zx1ua1wXoVMov0PPsEfCdF7Hn7rkWVUan9YatzCNsipdH
BLJtQ04b8cPEPRfJWA98uztXlUWLHgap7Dp21bG8WJGbxdkrm/rYo8mViQCFJlVrKD7v3cS7hFcf
9Om7Gq16KWT3Wkr3+HoFEDS20I/GJOFqmTDcsWZ4ba58uboHTi2plsguHxLNVPO8Mim1Stop/QiD
32Y2MLzJjP0fpYNXj3xbitGi79N3PNBEJmDP7RK22LApBk+ohYISihpQoLe8PAcCaBTHkDQ2C9yO
9diEh3e/H3x9GspLgn0S1oS3UdvZU0XbJndD+EfFaSOqHBpJhqSiRQrQTOuoJLoIMWyhXLb8bSgt
o2/TV1HWyXH+XEHw2OHlFB3VjrEHxTy7r1RO9MxvBJY8AjaZI5lY+CbMlTNMRtmE17dYzLP+xTsO
9r018UiJ385u9QebeiHmxVEyFtF4Q1XiAvVZP55pvksKiJWT7MpRxkVZ1yk7Uya5z8SPFVMC5B+7
nrhNSgKjl/X2VNjmwNSWLFjpwrRXfUX58XodDIfuNth6QhhdVsOBs96Kbw/ueH7kWT38faNM8PW3
+/KK/ES5VDeZAObdSGMw0y1iXny227jAV0zQET9MNOQbasKVkl1BBjS0Auq+PI3KB9bUQD0FMQqL
GVtsG4zkx1ta4jBej1IFMjb+QJdg/ZcIgGg0K2+M+9GHVPu9xmO81dzk49gTUE6zH2OvYcQufsRx
vWT90GWsE/60tueymapicl6k8t9X7ByPi/wh7A0AANQAuQ47+6KmgLHKkykEuiGFZJYchAdUQ0cL
TFikHK6svN+8Z92VbHxo+v3mGQvnG7P1ChCCLQxPS1UV+dvACe+48gTi6yYcitF3WTD+NwS3jDmg
cu9kfOLvSxdiuzVLvuQSNp4KWAExj/gBi23pEs13PsqUqvA8w0pUBJMzzbVnxgi98mmMGSxetbJc
p+RXvmQSQbMLNd1phKmJ4HmorRXI41QUr018D6BCd358Fn4m/R2FTfQpaZIM+m/np601ACm9zghH
8+LdIQw6nA/YuO4TxWSsq1lJecqp/NsM/su2mRv7cyFY1aDol/yOeG/V76ckqU3fgH84O9hvjzO3
Xgq3l6Ei1ENm0vDi8hfo9YcP+ZDJvnXkJislI5yrSB5yrzPEW+EZMrtanf2zW5HrnhvELku1vvrT
ojE+OtZNmFuxWpbJv5B953p5Ek37kbcqms5wfH/QfoS9rMXFVPA7ytWqpVfKiw/tqR/H7Mp+7AA6
FH91xqShVuNAdE1HShJ5bg2U4cdbA924Rni5G6H3ExG1iHmf653JcdGtlsitQ1185CfJXqcPIS/A
PeaEGLG3laQvoP5Fc3WOeS7BlpWReiA4hJipVOPN5ZbrpQKMjxYk5IfasUUgWHMcM+DdFsvjsj7V
/akZAvxj01BtCA/2/GMaV/BkZ4nZttp4Q0LIUxocnucj+MasiJmwFInbX9y8lSXFi745e7eqxaCN
gC64H/b3g2gkKATJ1PsXlEyoh/hNfiUu3SK1kPRosdVsBX7NtcfzyhPk143xMSTC9tLQvv0fsPi9
qqJg7hcVhpfP9ZA7BNWxuBc+t6oj0zb89XHOozfOgxZCAYcsHp8C4RsfqUArKbmo7gmq9EMYz1dK
RuljqiAsN3JpNY34ZqRBgTtBGYa0h7iJSBN3izpRnxxv3JkD1m4Mzua/2tV6aEKxlA4whMaTVHfw
a5IbShqj0BfOgEXGRHx1GJV/E9MfjavhcWsQX8v8v/FtAiz6EF2tmtYtRr2gtu5yxPvUcVJnh1TV
vahyvMbjzDWbkerpinWS8olRyS/jx7kOSPhQrZqrTgNQlmAq3hpdBMhXySKSw2m2G4/UqECwjfg+
dy4GTkFQDAhFHubabwbgnCdTOSTkhjwIFFULB2Hqc605BQVOoXWmN30huAywnvRT/eNyUQVPe2Ai
GxOtidx66azcGovFBydau9Bu0L72QMXZMN+EsXFCSiIAdLtaAsYpdl8KEE93szEjtPkpTImuKTYx
XfIruM4NYYikXYutFuCu2l+O1Ad5x0FHzxIxkYuUEIhSsazVeA2ypol+8S+PyXnf4gFtZFpgbO4+
0Gc3UflN6VySKCUMzUzMkoWGDD72pD3qPlHH9jW762Gw2hlQt1uSC6iew7tF/Gfan2KmzfNZatMV
KFPzxZK0XYZVpSCRsirQYr2FHZ0IielUThSYPXfl6dlqYzlvD+hkiJGQIaN7DkTnvhTQiQ5Ezrvq
MPKN+VIPI7RpkqU7pk2xLVZ1F9GUOq8LA8c6xxi4gD5eQ4eiRuGFVk92nwg4SFYb9/+FUgvCM/LV
LuzaMllZ2acjc+Bt8+m1FwYk9trKoioHKqKo4yAvocwAbDC8vVXaPjfPPm+nqOFILqS6tp6+iX+5
4DBVcyXfHDGfJjfqeURIVZiJUR/G1n9GGEFjb84oxZXry0MHOcKOi0XQiJ0R+CK1+XTAcN+EU4m5
6TSHpJvMmAzI8lfu0DFv1ySxza48iJ85fYmTSr99eFEv0pMWLQPqA9e/nUkfEXyzN9CaW+x/pVvW
Fk+LpFM9uNIr3No7YUDKXdpyXLoubzeUN+MjCSmUHovEr7on37j6NYe3nFJSHpCaGhi9Td1dAtml
BmAt+HxwktnFpwRGUUyFVWGIq+sipORMqVl3SDvGIxCyn5VOgvTzYIb1h1RkAEzU/sWygkoQptWF
aoGl7SEzYAdc5n/8HG7/ZqMhe6CYqiQF7d7iFUSAMcddafq1grQNrV0kUa5AuF01ED8DV5aZnMXs
3/BmRyj6p4LIKNpNzEXNe0obkQ/LLBUb3e2/4A4QBzGFVqCd50DYRlisePpYXtuV3tBhwmenMvqX
rcLj7tTo3jdUFKXhIOvBeo3iyqEtnhGoU6K8AfM9PFKAMV4veL5h7syAG8/Yw83Y0DxFjTHd7ylk
bhF0EqGK4owbE1qrevYTUbI1qRVnfoJ7U4ydl6cgXbaOP8S8r2HDuFJYJ6KjZJ4N1Epp92RF3efF
maB1c5UBQ8HKUy+eK8uZR2A47hMZZ6C0+6Wi6fwUBY1YoDvHEV/m2YVBCU3QoT/UFSiZ3iMeEhAC
jNjsKFerfdPtN0FwZQNUN+a4nkYXkpMGDSiNuHhI78Vr0kfAZRqHtq4vqsXvEE0nPDeqOXSkVPUc
leXSfh07uHnRkGmjl3atevGtKXhG6Llkn+3B9LNHjvtjjMm2/ehFcfXDFU252uXlrlusc+VaqFqf
ScVbrZxeWDFyql+jH/v8fgLGV+t1/8AFkLEV6zBSv2cgGWWrEQ6xmYeJDu8Px3Z00v4R9B7gXYzH
zuQ5vRP9zhBXJDVsOGHm9NUJ9LggA1Ivfx5RiGTK99VyelApgx0vN/tDe2N1J9ZQVx9UgSiZCzDB
wepmcn2ZjrCdGhf1ZjAbPz97h65Wxwr7tGE/runsTuV/G1gZI3uE6yxR7XYnHGXWfq+5p7Co0PM2
p6zPggCilTD5LHfI13TVX/IiLae6a2OEaJGkLmvOQUhrLv3Yb97svXlpFv4upoqwBRS29/Gd+Ja/
Jop4jMnOvVyqBc9VwFJbsNJLW2Mdm/KM9k+D/9WpIHC4pjvgYAoIJqgrS9yMM5L/A6e7LAgY7HwW
jp4siouUYuAx+6mLVj3lhlC2Pzayer106kQpZReazvSxUzRCLhQhnkN0uequbf+s74CQOZAyyFTA
w3aewl9jQOVBC3h26yf80QFcHLH99Sc8657REI8ysZ4cugTISgUjX6VtHGOLhBxpfX7ty1OiMA9S
YMjSpajHiPwxNrQbnzm4xEKDfoUFQgoF5sy9drx29aPto0g+ficURyzj93FULNlkdT9AZAxRP7rr
3moOuS7ig2Fu/i2TwcF4JEk7Scq9MMei+ArK5p+V5Ul7vUY+mnIm2iPTrVJPt5SA1JGkOg/LG5kQ
CHFO6Z+Jw0dQ5I4mlsxvcbyhWgNWRkFB8Vjplb0cH5Qfm2eMfjhp2O2+YL8eUfyMN10XfhYfNPFt
AroF+dgWKrLBOU09DRVgJB+eb4zp0fer65i+SpUQIHD7oXBDrYz4IN1bV3M1/um9uzAdtP5p1hxq
FQsNn36HkyA6kUpnKy5m5gFdu2BEQxL3JovGgOQw/DjF7oAnjqEmnYeuVLyq3ssHGZOgsvpc2Ylm
0Rxd6NgTmCxpgIX3II4WhJRLoLXanGZtA5fQn6QXgRnHXxqBi0BK52JBg4fWi0UnstpU+nvCt8fD
3zeWrQ5lVqxmKlJChyGdb+NIUrCCx9RnHDdJFoQymTkKrIiyg60cE/fUESB//J3WmiR+IftEIMwz
BlZ0sYW8PoI2wEPv4aqaUEnTPmSAL/u9FTrFnqZkf6Bz2UcFa9TMELoR4YddVTX+jWybRs7bftL2
cdVlSnu05SJxqW5wTt6H4BqT22f3DCDUgvChVitXTFZdQAYTJr7ZLlFL7DrV+qzVyxwqSQjTl2QE
/KxPWHFkY2MNoRklbgOhRgxyN7dkkEmclq0l7P51qBbjfaJKxbPhm41fJphSFerkbx+3YVPP8yEj
HIJEZHgMOdyukjt8YVleg9WdWKsGwI1TyUVv8WtS3P9KkVdxgYy5j+RCovwP8qOpNhR0muft8Pq3
hvLn2Yjcfl92wRQrhu1ixuYEvcLHhU8se8dokrk93ZBDQ8COpNJ9Hs7rqtlU5m6Hp8dQczikDcvL
M5HFhnq68PxpWCJq/7+bSzt5qb2doOCgey4xKOe5pUJ051YIMtMcKNsvxWlns25wWR/jeDGy1/DW
ClVg/g5ujHhaw5L0hyzsQR6mEwv3RDhh2VBJVlcO/0KaNmxLapWqz3XCYD5vDusPtqcBNjoJjLhG
TywdMrxAceRC6O1xPDW6oa1zkG1aOCM/0a7fVq7Sdz3qhKlMsSFyY6adp8s38qqqBQiwBp7iyMVV
aT9XDytpqEObgJt3cocqauBPjpe6Wz0y5D1GUR1gjgf2NQjAOU0kht25ZC7IFAZbPX9cI3k3/IL5
xdvVQ+UAg0U6VF5s3ChtVnauVk818ZVgNkps+VSqYLtNUcyiwnPu9k+x6OBJHZ0UBGMTHtd42FJU
SZ5uD/S64ENBraAryVUtNVjO1Eb9lfohszxWZsmF7BSMtvv2YQkdjvc5kRAPuueuleJnVN3t09n9
Y8PMS45+dB4GP7eFZPLHDgo9ahckUX/5gxTX0A7fCSNMfNiaW6pAt0Mffi2hCd9rRER60u1pXIyi
flO9wRyGCZjoMhqa9iXzFJanbIB2hfJwFH84rXf42xlh+WCFm3iJs2BRb+p4wfWlQGwcMEbsVfaB
KgS3mYS4enVXs//AXF/fO4ye98WFN+M+XHYPObqzen0wkQM0Oy6Hy7Ir98WmWo2C8Re3RmuvyAaj
Lq1I1Y5Rq0tHcWAeHhp0VIt9Z9XrWlAjnpLIwtDM5MSYClYwdLt02gu9I7U0/IsFa+F88XZxdxch
97O+sKCENg2D8BiGbKxUYfY2DyeubNfFx7kBaW9iTFJxU59P8Fheuf2swFBUgbku8QELZ64tLEjA
4AF6gQ92a9KQXMAGE2p70TF4CkH5GNS6iggJGFvcbRF8Eo7FXpan8f7EUqJyXUObpI/1uJY5Wy+t
OVZxX8Reou/WN3LRIrND5vHDsjSumKQQfcBC5TKQiA7yWmURHiy27PwsCRJHzNO7OLCSfSxV8nu+
JgCA62aJKuPi2XdON4j6ia6AQ5q+XQQzSu8adlEZh/AVuqUXQtD5sgKB71Z+2WahwE5P1FXrG+Km
gg1toVpUDEWZ+mtghHFug/ogxpKmDkQadwK0q5rfvhSh753hf9cEl4ZdN3gFrz5ZG4anvNMLlPPH
vY32LCQ6yUiIZ02tb1Uax6RAG7eTv9iEXj22A4UUwhbmz3wRtMXbzm4mHua5ESGw+rCVYNuxE9cI
kIYp0/gCXKxBg+KS1PW7R6fUggFr/KqT/Ef1QpgZS1TKkVQQ6Pu0xBa+HM/e01TXh3Pc5U1f7XjB
6pS5mx+G1Xj8gi13nSR9sdRNkx/jJtZdAOQf8NGgxjNk7q8O3NJeZRtCPIK+Pl7+TJ9oBQIUDC5Q
W/T00c1eV+xuTPy0hlRJwurlwpG7NhlClFEhkKIPKsBMYEY+yY7yOOIWKK0Nq5Vvd5TXFyI/2N7T
l25vxhyb8gi7hClCwYS9pb84XLPBY8E1MsoHl7F8juvolwaag80jZIU5HobQ6fmgZ+wxkpTX+s+r
BLm24tHWx/Ga76vo6TYrhj7N6C/Pj0oQufSbWXZcJFh0z9sITl/z3zNtCX6MI740ctVaLBYPNEmg
vOWpfYY+/nxxninCwn8ZP0nZvW+xXuQalEKPmrwd4o6cTpcIP/+1Qv8/wzyIYTTN9S+rpckIDHdw
/o1df4iArs8m9B1qd9ghvGpzLfsE5zUl8ex+f+MPFz3zKByDyTdaYNSQ69XRub9JSW3/8YXFGkx+
/msZZ9FEIXLHqmp0nk9os2kfjYAPYQaWOPIjQMz0sbgitrrv5dyZngUTBA0Z39wFq1anpD+VUF8r
iq2ven99YeBkdFY17EPtCEP/J9zOrYLGaUZuCIzbdDpCF8AtUh71IkcMG9vWWkVDYQ+2deKfMAMv
TJowzpRUyhZfY7LFnEF7yvWTR9tktgssSjWp+iViM3nc+Bk5FzUcpEP8h5xknEoAElZVenzYI71u
0bW3p2gy0MSon1i1hQbwkWQaEJkABga1fJS2hc7oWZUhAKtpt+XHJaeSqCVobAqV7PstLTPm3Z7h
bokzlOMbzjSf0OpRxRK0CxDeh9GRJHAMm1/NPlOyMQtdGvGYHKOQKSh7bvto0keKMpDlIX1vYSK0
ho+mKmu5aLy7IsTZppb7eCXbVJ3o6EvlC/ifATAu9Ku3H3oUSc0grJZCuafGE8qBbgHxzYt1fh9X
/3/w7GrrnNzhOY7XZ0GzGpbxoJH03NFuoCoFrl3Q7SDxjXghMidvpacIxnBDofRjqiEbrG+9GWoa
`protect end_protected
