-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
H39x8Q+zyD6tnjVV3voNfVhNOAfi93UG5uMsGC8L8hIqzv4sfO8ipqFwBQJUItkJSWcF4yQI3qsz
CZbvtw5gCS3ROwgqKkvxR2ag68pYsyxLfjwJWtrbNKFxVOp7L9PGrO0jvIv6R2cIUBPjbiyDrPhs
5x56LZICgy+kab4lrx+ZAqKa1ms8aPvN0hiKD1mYiVwXNzk/0sLGlq6buayHsa9tJV+2xB+D4o9A
zHO7Xwu8s9VcigOPgXJa/oKqO30KlOAX0quBUWVnWvlpvtJQfXIaEP/vRaMub42/QzWLJJMGur0o
qqGDLPvs4yGhR/k/VgoH2yvzYK6fvwEhbjg00Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1728)
`protect data_block
vT6D7R3xan88M4WYoDOVGXRWXwuo7z/IxqZigFPwLhi60qHQbHsMULdjqnuMol9RBA0ZyjVyHRcu
uLEbukurJdPq/t+RxfC5h3hnB2yodTG1VOFpZBQT1z4VN/Q34fsyFQUJxSLWcFMaMyI0N5jbOm5S
Wc3H3n0mLJ8cr4F00Q/z5yIKz/u8YiuFM+GhMumnlu73+/9/a8r3/kbqKTk4+F0rMB4NFAe49Gm8
BObZFbeL5nJa3llM38TbY+fzH7BpH3wiK9HH+oDi6RVKCNMPw+IjfdpNFQWmMERam5LytvPEiw6o
+1rrokG/e9R23YBS32ILy1zoDyWVs1exFdCD5BXuiKo+ADBXeCUrfllbiQWvKdLEgv1GMIeL6RiO
BBDapz0sZLSymXlqtU9N1VAVtkq7qLXOryYbmGpNmZvzhaLeBk6tqhf90F3CL9Z1NXvOS03T9Tye
+fKg74iEoiWXJgYx08k8P7fOEk4rCSqCAs+09KiyWru8Hz5PpnEXivkkBV1oQXiJ9hwFLRhz6jgO
gVJPrE33j2LN0NYmJpVyM73pU7hoEgJt7TcB+fOKz/CvWyBOcD542uZ1LBLza0iSUsrmwPALL9je
zqHwRQFlwctXiCSPWt1VYhbDOqOSGQTwsYBt31FJQpwRB66M54ZTKUe8teP/eEmkZuzl3nciM3zr
zvlErO9Ero+cTdzn2QuWMtCXI2/+oB5TH9V7naz+2Qfqbjlm3zjGuzSy6Xpma1cn8nrlO1o0YgGI
qARJGXI8yrJnNW8qBXEN+pabTLJCYo4R/qoxxb4XpMwMZpCbflrMTv7OmEoLiBAjTGazjsioOS5J
obPkJzFIk8wgXF078cKlVeFDpI+oVNgGo1MVkUSAEh81/tUeYKzTOt1CBcTo0L2zE8LajycVyCAN
1fzgamB3olf8JH2Q451mEoOtXwroUy5W2UO5cq5653g1CWttjaKsbg6YBdVdWXHb8WDhBIWfmWyC
rs9f+gL/IspJuOCXeygaYQeJkFFj0scuJs1g6RDh0xvg0EB674nrfE8kytANhcnyvLYVJeHAnZPj
pI4h2j+o+QBlhQQuowRoXWS2T2BscQHo2jWukixGE57YLT6WlSRj+h0TvbzjC1Eos5w0jyzf+69/
vzlpEAHlFKykTCmXhxSJUvasKKxN+w74FK7RTbNZdkCDmgH7Yrzmjmw49+7eWpDMKEGaHJJt9H4Z
ySr7FusJncuAh7cAnMoG4JNTJ2vzRpAYGfqyOnzTpelU/7OzgBSArLnNqggQ/V3xUl3mdXdxiuc7
PdyX+slNEbGd/e2zB1ceeSB6XZ1qoDHHti72B7iEgRqAFZhxKBLOwata+EPfSJlGsRfQ1NAAGmvI
UE++A4IKu+3awyANvIlCG8IuDPoexjCl76aLwte+wEzpx5EslQ21uPDVJX3HR4tHPZVwvhg4DSki
1CKFI2G08Zi/v26JrT8pMjldmpetRahl2246W821pDBKPI3TC6Ag00rVI0hHB87Tt4LteE6Ntark
D8n1j3HnXhxrT+tLlD8mXDpqfxKHREp9jyTc7ltf0TVvBnBTVmXtOyAqUo7qppub6OFjx72cYPcZ
Lg5c7f5aOgGW/OEdHITGzkY4E6vAMUV1itpYJetQdijlPxDS9AckVweN5T1A8qG9tS7LjSgWBK15
K2GuZZ6wQvSN/789Q7JSNzZRtgLUkUi+s6DjQeH4/nCIHDKWA1lydJeRwEGkIsOBwXbU4b7xi1EK
iHJxoftK6zvQoUplW8dDGXrIADc1zegaf2eqAnmiBgpI6H2hGnmtpwu6j0Lj2hho4/xpfzzKZRH2
BHIXmLmSFuiie849m0o+nPKzQhY6SpWR/kGlfIGtGfVlj5snZpALuGP4L8aVrCLoumZG2BmXrtk/
RG1eFW6s29UTCG4a5UPr7By5Mgav0kVUmv55aoCHkya0Qs8WOCChdxGGR8fUwtX8tWQJezHkJaA6
SsZPPGy5PclZ9KjzI8aM/DB7OA69I1bLpOJrlmAZIWaJAYTxgZRwTHK++zEvdi4dD8B21EEPPhhA
luAhSNHqErbaNBlp0xRO9ieC/74KalBeX1c3sDGOE5ybkYdYUbnACcTHK/TDNkNaM+uZAPI/vD6x
QjZ8fVyeAPp3bAKBAUrsvbuzdXsDq8yom7UCBDyyrwq3eC3bMmZRz6uKuJ3dgpTevYNw00uIWjoQ
3Vt5eOLPqiCEstDSaayGloSOa5jdtxuXGHJI/BJBg3lTvMUX3ag5X3c+oCzk6GNrDmatQJqoHosg
c7xrICmv4P5Gi+BGL3F5Xn9D
`protect end_protected
