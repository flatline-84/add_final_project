-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HRo0f6jcKrFHc/lPgnv7H7PlUGjJZAapX1XbKjSLWvPpMIeo/+BVx+E7+HpxRK1DIAq07mvJNbG6
6mECkhCurBZvH+cfxo5YsNB4cNu/pSCjSv/fi7DaJpqDHOgHrEi2Yj8m7J0vjSptIwvn/qwOaFGG
Uan1FAm4HXVd+JGLcOyP5vBrLGFHLsLjMNaIqLeW4wacVvANFY2+6B5P/0izaCMm+Y51lTATHZHD
FXI6yf1xtihxISFpsE6ChxnqiAa2NeOxrLpQ6F8R5LMXvvllgjc4d6PIsxQXRW7r2jWYpHSFsKW/
b49Ca4j7f4KCuuiq/wdorQSpI4IDFVz7FrEKYA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13456)
`protect data_block
9qdh2ZN/x0Wjik9qmh/fKhDEmqWBsPjkJh3FZ0qHMnpU4cJBWzl4b5/LRZ5Cjud8kdqTCXOmpen8
hxvXalFJze4Jx7H8wL/wWOrUUOWoqv2vpIXiHzHyVEXJ6MF5MZJclpApVnkL9qc/IS7CXMHbPk3j
fFNxsYss0CwSjY+Y99dV48B+F7QqWZK8AOErMVBet3KjD7p4dc1Oi1cTyZrUaj2U4+QKcWzM0TEX
Fo0a/0r3DEbMutlsXgkLzHlhJ8YrkkOWKxHzpbD3D2H4BtCXwte0vE1ZGx3vwvzOGGxJfItEslSH
sPdp6q691VUWz+s8mIt67sY1ZLaLVzXXrY1ZL+ZL2OzWfaQzrfJXDLRTSj6Dg3UwpwD+EkuFexBG
JVQbi0SWSB9PoxHgEYMQtLVfmCKCwDXUhB2ftkaR72QxYBEjU2DEs/cM7rJ49tWGmGZpWRRr0Zs1
fr1N1duy/kBTC0ILme9a9JzHxpExO61fe/CtseUECkFtWQpSbdkMfnr5EbTOXmAjuTZZeVICyLy/
ozkdjXLnCDO+BZNGU0clxLnNYUYn2y5Hsd73M+fdL2EOtm4IyNxcwUg2p1wNEh47pgNRMDeHTCzw
BcDdnANNgCHDOYDIFpG6Hg19KVa+gv6il490mSz9ChQgPP0/qEcA5hiKf++pW3oECc7xlnMQ3sBf
SScYd/bXNU+GLU4frSlZp787h+hOFHEGh4OsMv/gQScoQwKwM50tHyQHkSmgAi9CjXJ/q84H2KbJ
NA1Sj6Cry4EI0CSKo22OcIuCfYWUgr8t2gQUiXoRF15uu1OVghQqxQdIg++ZxnsEkEm5JIugV6be
Bt+Vi9SHNg0Cq6qGDMKhEj+h6Zk5RzHgZ9lwQPIm7rcgo3Zem90pDdNgPNj4ThmlhJIwUBbx39ZV
nlyk8L534E4RiZTAXrYfiLt+kjwJFRgJrlBwfjqGNsDe0cG2HNWWvNc+733yBYzdQ8H6QyKqPyfG
GFRdVd6LIM9f6TmrXrbcQfDOZHOa8ITtZEMvrRBQ37s4uyRXPUGYtS4DxwoNGY+qoQVE9TEIReXg
VTwNxOrp41IkHy5WDT6FHBbafDTfJudkCos47t7alA6WkuD00nxnJUOEa3FEQKXKKHhXdmnfsFzR
t60XX+Rk04zLU+IKtiQ4oQDbNCimw/DVrGUrKc7XB4jObRP9uFMQ0ZkOWY0CQZ4jc2w67KOKu3K6
HitaN914cvOXeME81SzQ2YfxNzLCE3gO1tRhDB89+yla0CMHVFZ5scyWWHpMfZK5axri3vXk5soU
KA5gEydPtzCYb7nTmrIPWX5yfsYveoAT+ZEu5P4PS09VWh3sqAkeLnXuN92Kt4xbyKGXizLatsGT
dR4KKFwUCJ6OQ6be04h8hPJjfWvIK+PTu+xG5e1nWeEu4vU2kuPwE8UiDTTimySHU4H4/gdhh8hH
tutZVIdgqQt8cm6+/2HvyqD8a8+QYR9IlCRSKC8lckYvLPCdUpJgQdibc6tikQ57jsyNM7PR1cWq
76GvGkHQ1UV/qeGVTz8PJ1/uZQ5B6iRMxsj6/1al2W9JpuYevQfH5OxAdq6pR2JfF38xbwQAXaj1
CmexO4uOYlcEoIA4DCHeHeyZ5mnn2c7haJ9IrxhZ1jIP1Hk2nV/w0jevM23apOH2ez8O38GZsHs/
w7yFgY66tY6iIsI+kw8l+jLhLZmHoaDTuT89un0Z8+Zujcsg81vloTmRryBJPJYRF3yjnYhB4cDz
xTkeOHC+Pi0m0yXypWUl/2oakucPV3sqNBM9eTt0G5rBvUD07e5MVbccUTwTD3M4SV1QhQNSrinx
pfC4SwplxUhjGK5Awheg5eQcObLg6bVVX9EkQW6ur12YXeDTjHx3d3sWsy3FFXwlvTWwFW3LtTsw
GDWnj9tPQI7wH/w22Pf69eFrhXddRfm2ejjxmbqO8KiIOoEvx8LQTjDSDR4CQZnzqNSk8NKtnAzJ
6c8GqdTnCRU0K6fo9zkqO8CkmbTuPDtWKAHn2coDXbL4L//xnc2sUeZY2qe1lyoaSFEFE4X3fv/c
l7DQOJh8XdruNbaxm98sPZNSnpwaqCP661oq//DF8JOB/UFPKSGNKlZaAIHCYF7lV6kjM6TYqw49
J1lupgaaI9FiiiTo/W6v/k+kX2wFaHlaNeRQU1ZTEmCejhi49zHr1U49t5OkmIcO66sCzoGWI5zD
p6XKFNxN5g4Xkoy/sHNxUfwm/8p20MBTbr8Mc5c5/CHi+qiIzXlJD8AIlydaTg62K4ioIbk1yfVd
tVZXMhwWUYWE9jedotBoZ7I/2pG+rxB8ucR46a+J7UTlIqTj8chMvo8bxJdmXT4Zjp4Tvoj/Eoc4
TMIY8upQ31pi8L+PveOtNorBJNyutHPp397xS2iih/rMGJFoXn84Ufzn1r6h4af7u4qRYJYeAcTf
rXbBYCplJ2Us171J2xPvRRXzZM545Ec+ONoGt2V1iVJp4cZyAe2oIvEwHTU1LAr5d6MnupICwLaY
FD8161lpv1OrzHeGGNCxg3xmhtQIhPCQx6kyBnjNnwJf/uy9Bqb81SfrOMI8p3hYC+qhDPYDRGtw
LP9BuGCyZfFSn8P3BUzRRRxegs896qO6gw1RJHHquNCJqS8A0pDS65uhiTYc3ltSc0c4KmfolwPO
VFrpMjzS6UXPCqEaoY4cA9crYzZRbZzZrljsMon5inqss33GcKwV+dLUnkbur3L7WWgBqZmCgMdt
tZ43cAQSEIidCjCQe+6BoUhuJDjyW/AtSigXK9TAf1ns4Jsxd+WWCzLmwO/YapsC5tWnx7qwyU6d
Qki8vTPGB0LFQoEDZxQ24GwtU1QK05X2+gdiRZ2tyXsC7UkV9qKTTGk73rM5M/McD8UBpl9PifZs
Dtei8Gb0RedySISmicr3De2mw6Ujvp7xYmXpuGSoGfJ41QIHWeJBZiATXrBFWT+HdNNlQZgwrzJX
xSxdyymsve/2qBPBYRUcZ0asYz+OQmovqPR+B80n3WYer7q4q3E/Gk4CUjf7dVkAIA6ImZaWY25q
kVIozKNLqe48rvK4pXAELY3YRLtce5iwi0j18hFgdhUKtoIK8qxoZjQC5LVqYnK7x5shPq83h2K2
ZmL1xh9he1VvBBVz68P1VuFkouXJ57WFiIEz+Pz6w5z2q6OGTbySe0R3qSsO3BbxXZA09ntBAID7
BK89RePjukC1GoYEOItmpjZkkiQTyqy4/iJ7pFQaKGGRViiOx4xWKum7fNM0np6GTB7wt7yQCNUk
VriGCgfpIVRJ3m95rJORwsNzIDTfp8itd+RXX4ap6qdRwk6fUZd/1l35vFjxnt4pP+kDULtjDFvF
sm4zMADGszV9UCk80GlaNgQOPh5yI1E4OhOMa7US8RaRS5u2zel3GopnEDdw6j2gdVDRJgDjzYZJ
bwzMarS3Qe58PuG8sgD7ESvWgUSKc9AJ2kNOd98hHJ8eBiu6jl0lFUAp7YrC9iqEgzgfGpBYazW8
BK/qj1uyA8m2ekfav2WLZ2vrklcBiwCG4cgmUwEPMfV2uAPkbl5SxfwHfO8GfnEIS2ABnXYnvFk8
EUd4fMILATHF6aDoXwEvJIKLYw/iiCK0nQKBDZ/cBrV+hOBw2R2pfAavnHAu3bMThr0ojR19kbee
s5w71X1F73t1+XkFdNIYu4N18gIH35PeMghZ2DixpKvlt8mot10lCQscWQ2CwY2ZXp00Mf3HumXi
DOsaTXhjNQX/pBlQLZVwAxYZ3bZB0d8b7Yj9xW0l3Oe2uZUJtNaDB7m8qEBX8Fmw9mhzS3QYhnqx
Lms1kS9aLLN07ijU+nVOygrez/4uJAR1RHseX5F3CZ2Bt56LO5U7M/HQSnbNcZ5hOSwojIIryEyq
ZLtGUcWndSO4QC4XssasZyepltlH4lvhdlbHgD9ujG0nKWXKHrJvkcY9+GWbMYaQBZxQoh/G6VuU
+5YwnkNNpsGOPRvYGlzHNDkb9OsF1PPmbTxi5lrCekC9bdttlBWWQcBV2DKXh7ZMpH4v/KOcM9z9
PHqLdN7M0sJlkZA8JG/NGdw9F9mA/hcrupnTNDBc8oUgePNp+IyKzSK0wDXU0PulrRYuKNS5jnk9
hDECLLbAc90vuupFtJFEsV0x7SG4REanu7naQPXMzVVxF32IHploxPRlmPSIayXDsnbU9jnH94Ed
tJWJtqREp4Tkb011F6+8WaFUfRFJ8NtSOchdCV9r7MiH6SMvV85v2J8AHI+IiT6Tae50vpNecM1/
6FFFZjAC1Qtu26seHSomL4GOBxnbqlOa+OP12tpjdKtTSWWuJwttSmIM3cPHqcSNIfpvgInKw4AM
9jZhf3yWEB1EabEIZNFEgWsvw7H6TLYoMzvC6rfBQWafT1X7PdxH95XkztsFaMNZoG5gn0w6tIFe
AyBvF2r3589ETi8q86n4932RSPMmATtD5T/cFVfmGOZ3sxPNEQb6vTgOjmn93P3d8xsR63JLtVHZ
wxxNoNPetqvtxVYYX4wglVmdPE5bElmH5fHvQb2u27O2e+mg2eukdeJFg7T8aaQYdBKlPUq4s4PA
4WSBTkNjpQLw4iAF14RzRBqNsuAj/oKb21T/qdWtEKODexzTz41Zt86az9hUh43eGgK8cqNaO3hB
A8i6VRxDZJJzAU/eEVm2uqggxhhrY6GXVwufjSphbQaJb4/Wq039+/D+nN/9BwjDyo/u0Cf0B/ZH
zxLBOxb+53GX5GJZJQiEkGdDXGwPmBgfPdDXUysrixaQIyflQp5Memx5HQwp3QTDv2D1u2arVkc/
pAeOaav6IgQjnc+HzEa9oufBFVN72mly1u5OpB2c52HMc+6i8pg1SrH3fDpT6drOP4Z7kcb0iLxn
gWC4zNn42IK6yPLIJd4wOiYFpSmg/Wb12SSDJGLAaLPjCe8t1S7RE7iAunjya27sYj59hdxf36zc
BdmNxzP3YgsOpde7c9fAp7/Petoub9v3yrwbngPwn6faRa65xuQJJhn3HyjxDFmfepeL5lBIfa9H
GDXnB15R00kcyd+FJhgUQvfdeS9BkKi7TLe6TfPhRwvmhpd1/C8i2qa7H0q2pIDG96GOS/whqzy0
76KvidTFo38sqihGZHU/+ZbmQVxZt9cOkzm77DPKA5aOOm3+EEjRNJ3fI0i3uxqJvpAiVMi/Wf/G
PM4VGvMoKl31Gz4tHQgAiNBqxRYYsRdE4WAsbKpF8CZoAcpMzhaPTFsFCga4+BubH9dMvvfaMfig
vgLQMlWhpgaTOewVcVlnvRjAf3vGnCEUpJPKbaqC0XgAJr3eDBb3UdnPTk+7DzzqK2BC8fUmjlt5
8b3Nqc0f5XhXy5/uM8OPUIND7mJiTLMnTWSdmwlsggQotdtSncF9gCHliRgVaXN/fWCVdgFU8dSD
G71Hg62EoOo0gcrehUdg3tNvewQNZpo0naTXAE4VsEFpRrq68pR0rh/XZ96yD7EkYb1p+UXnhz/h
6aF3bYKjXXfV7slWga/okJ2Xv0m1ZTUId50td6tQ2hMx0BQk5XB+AVmOlrEARv8yqymMVYJ6sEyZ
paiLJvTqynNipBKuPEXixbjRHVdtwNBfTlKwSjQpC0zFwbb0RYeVy3jaqyz0fdMnfTOTACsNzWQi
llQSXAPbq9qI0VEWggXL2x9AJWA6ToFXspGX/ka1l3glzdfGgVXBaw4/OvrsFJc1YMmZh/sEJrsR
1JOgNYHlh2twSLtoOVOhjfaRFbNIRMpX+2dFpdxT7TBi4Bw+zPpA3Yt3FK7aK3Q943/aPrBwX0h6
v4EO9ULtMHhtGmmPfD24byr1//GIZAggoWWRjeUKt8bCK8MmraBf8NhhsANuiq1QACkiENDnXo8q
I7beAlHlgxmzcHOHTeGwpUZo8k/kvrB1oMJjeQtDV7NHBrk3/9KJmk9T0FXvQAmwUePBneqbqTm1
T/sbyCNUROtr/YKY1d7v4uuEIbhffbJds6HDxs5HX9h6WHgGSew1UNkvTxo4yXJwNNNt/U01OGEg
oEM8rJqJTeQyckwPRz36w8BUWgbpIqY3dw3wW24QIrIIczEVT4ZHj2HBGJ6wWes224xccSHaG9pV
XsgNX554XV4XdQDK4BrqmYj0mbmcThHrrrM5kdBmIHBxH0nFRlB+Si2DanmgK5y7qfnD21a2aWHX
fOe+TRAO/9o6Qk+FMpJISmaWIEeb9avToZojKYxtjLqcV9D2KKeObfg5p/VadIRg7CLaZyD0aU1R
pWGi8D7qdZ6TZFcYdjEw1fvkt4dP1yuCmhUyU1pBkLlQkT1MuPtw0cYAgptcjXmoM/JNvloVi5xO
c4aVigcQ2Vl2B45SG9UL6xJDEgb/VHDge0KHDqsZimVU2mLQX0cpW0r2MGAA2a1+LMqtdbMyEfkz
YrzuEqGXt8N8lxFDEVGgMGgEcLh3jWY6MnouIhITy3pVcISWOhwSMYZNpipiyAvhFtweEKk/ihv5
Bp5Rf0D/dM1WS0xigkyFIw5zl09nF496RvGy3bwyyXIgFuePcSYobAUJQeM5kqSCJJPRkWkMjeZq
u1AbZgcosRwtB1zTXz3bi1hzTNy/xxEI5SRSPej4qU/yhZCJqRyXp8ypKg37iP14OUwmGYISQRTC
SprzKFknW39H2hHjvMevNGZH3bSgGRnrMi93416mXAhdvAAfy0BQX8WZiMsrxBZSxOP+uICJ8ScE
EAMTkBdPP8zY2eYOl9zd2VX9amORwoIJGqZH5lNjy1/9hjeuRbn4iMAc7kYnPQxdo+k6H3GyEFng
PO/XbAcjbHP/scPp6KzOvtHGX+VDXcEeWwRyA4tP07vmfjIG8d/Xp50Gdm3LmD+Ryu9md+oOXEOA
XJajUuPixbE220F6BKojtQNRhf8IApfu/7q+LT7UmDK1r5FbAzVOotwMoY8NOugo8ujUYyFwSOE9
+u5/xqUZ9SGH0UzR1avr5T47kTtfjJMUqO2/sjKpYIh1ArrFVo9Z2ycxy2Mtp+7d6owDhTKOicEw
ZQL1Egmyn6zOJE1XTuuaqzL8s98t8kwjbDInmUuIrfQg3xAxOpyBFwZiheng/4SaSq0l5UsZa8Il
GVsc/Kli+o7THOA7XLaElG1/DcOc5ZVPuU6NM3PFupZ9Lz25WSaj82JN/5GSAg1taUIoYkgdzNAW
NKFekFwEG3rVplM2SprHRgB1fxT4dFQ+f5u/fatGbR/IZVyQGx6rs+STkvX/Cr5rU4TfUjPLEJl5
KcOD9unLjF+fTfr9NdKQH+RKjWqp4v4lflls0bdYWtBNhXPjxkJUpXitb1aUQTOEySRqZFFeey/+
4SaelGNnaThujWnR61RmajqPE0uxFRSwfJYcyrX+/e7ezEcIikVB01oL1usm/6RaDyPesStaQGi6
C750Q270k06lFhkpWDhHYubaEIBjG8CCcPszbYjBDM9j/4wUDgUqAH5Nithc0+sbupn9TuhueLvs
jCkiuYdFXvH82X5D68z4PIThuUX1qPQ7n9GlYoUSFr9Ef+uGTkN6uCfGj6tDtcKZX2hj5B39s7f0
3YMvKTDnlxEQM+nDdOkd0rHpvJvu2jmHYSTh1xg9xiq5nShSFh+5Mg05MbLcV5GGtuaparjMSauQ
FBpEqN9eRqgAr3NhfvuurxQ7qzpC7CaMGdj5t/xKk7ND7YMjHpe/ArX4/ipBSuqaxhZ6k2WIe1M3
cn79XtR827MHQBOUnq0YSoDTCK7fxwvTA18TdgHp+KQyuZRHRbTSsoRUP3j2jswen3pPBi/hHlkD
VzIQeS6cFitTsEraCh8MesM4iWzPq3TD0mGrrA11M4NLi3fXFgB3YKvI+6tD6vViF19T9gPB/UqO
WhSdW+Ar4UGgVnVL0RU7o3FW3oZJuiAyh3EzTim9WjOLmYNh/vI85hJksOTJfDH8qDxag18pXu/Z
JjB9/dstAIe/h71t5hTLdV7xuiLLdfjeT5UGysA0LWIK1Mi59b2sQHm/s8K/cFd4A5ld4XhnBatj
a8qkepoWC+lLdMUJautl8qrPJnIwUA2GxmXdgvTZT/pwDEJaXBFpm5sxJy/+iXi2DotHytjF9b6J
6GIpd4+VTLI6E7W/g+Cbgco2M3acBVKlpuAqItdAuHuG5Jox2wxUorGRafxPEh3kf+p5Qn3De7Lc
GcBhzTYz4S6bI8eN/ZZ/GhOyPWgBRe3MMqKLKrgAShpxesWuUPOYC9PBkAhkpBo35+gK8Lo4m4p5
B0CpULpkEwy7kteUGVFJPcOSr3dDyup9a+3F/9/LZU12dpEFMUPafNJKsdbfoiyswACB1KMW5N6+
s3b0PLgp8eIhsnsCN5yCxqqK74DhH5/sgiBeWsWkzEZkxmoGzZ2cCFhP8c/ooV1WfwJU43ZvdUsy
w1DEV96cKVmbR75D9liiyA9MJb/tR+zwh7Pflr/uiyn7RKdnbpMdsEStCF81jwHNxynEjpSZrNZ3
VjjPx8uDOvdxwuyh44X9jdVBmkDXlbR8U/F4/x1bf25loG7kAkPCrjZ2pvHKWjtvKyMl9ksnAmCZ
GQedNLMxoLXeMlj3Tw0toFJx+vdVud9+lDFn4bJldIfL+EZ4DXAa4Y6k5pyy8viOALbKkThUIHQ3
DanD3Ks4vxHdK6XGqhhbLnvwOnfZjJfgnH46LFvn33Ar2p+yFxSjhPrhExM65L0LDMXmPRgZ/Qz6
/CAVPGwcOA/yUjtLHqNFZYpjL7Imc72mu9fGmiod/y5ywMNGPyCa1JT9X+ZUmSOrVKq+kjE2lW5p
bFGT7fFpcTAqo8ZWzjR1OCeXexOF5JX4sBmPZKtZHFdNFaCXUGhG69+YOOWAZ/GlIiQyO8p9jn3W
Z6+K1Zk9bisEAPT8I+5al7BgicZogMAK8ZsAapu+FoDB0j2R1VwVdfd9F4NkefkrVPhk0U6oyiLu
DtPd9moyE22A0jhv0vT/vuJElsDzNTpK/NZrB8s9hO8RcYnwTkYSyyLMdsV8q+DFI2mhAKkc1fkY
iHK9msjPmTJ89AQoZc34M/q+y9kL4riRskw6KLkea0DKoknEzfRXLUUQpCfGQ3LBvrV2E1B2MGZx
HGzbbl8XIVNdyWKiSPY+Db0z0wJhVrRQfmWnp5ruQRRxx08gIdI95zPmr8Pk9GWDFx1rwnPcQGfG
Jtpxjov/XxJtEdhy+kDijivPm4HRTBKaGSPPILp4W5MgjOBa/gQNPRjPWylp+/eogu726QzlREz9
m/NjBGqxuBgCUMXxrgxQO9ZdH2nyOy2qOFkoNaoMNl/HN1YtFyLY2MAo32bHp3sCUfZqoyvWcCmV
BpjlFQszYvbgD4zoMdneJx7Za4KuZSfc/PTWO0gr0HEFYKI6CN15DbBTISIRzYBkNOB2xsbIBOus
kI4idR8QnNgF04XmLSlziK5zJiUavFmvI90JdP2AcdzYO9ZYVLH9/uo+3KRVZhjJlgdR+1iOaTIi
aEg2/0tXtm0gHSYc7UY3k9LG1wHEgr7YB+KurRviHTqwrSmeSiA2nMYgzZgopCANk9RNK34cS0c3
V8gicTg+FF3uYkJIMS2BMRsUBnA0b0lP2QEBTt73LUdWYIOmNq7/CE44lAb2bI3AciPJTVGNTNlj
rghsJNmBqNWBrslx8kLBcc8ce+xRGIfDwqziN/Isip4NOrN1SeB3jacCA5IolXKhD/ZsJlveYC8N
2smqx68JF4XM6Amell9eeJo3vRnlL7ZVFKq4/5MvcaXFfeDVUF6Xv0lLX3sSK8NaoJVkS0+O2Ngy
3H46Dhu9I0JuqVDUjXLIKwilJfpZNX+XGNTI03eHPWEDgwvPNYyavjOuCdtBSA+WEqcq12GUFROT
fiWiWX+mLYMq1KIteYWm6nHwcMF70OBXfo+QNKJf6EtvN96plJytCALA0yafRxBH13Li/vM+dgRD
d/iVxUqC1S6pmbkcMwBt7Ov7lXoep+FiKmMjHhYQWpChVU9v/1gPh51t8CT6S7pgS+v+9uj+JA/7
Mg6Auk3mWfZMeVePXRBsxuQ3JFWi3XCMEQLDGzIoWabW2Ew1Zdrr8+YT3SrKDYHZO+R6f+XX2xJ/
LpTVDJ2dU4uB1q1QtMPqtgtfLYPrZmVvnfrotg+Nt6fqljkTzupo+aHhoIRn9z1DSoDqv4oo7oNB
p+HZfE1FUVySWk2VHvwy9Ov8qy8i99IFxgJKJUjvNKT3REKLvljloqDnS3NqpA+jmWnlT5ww6b3R
GdPbK/ko94rwaSfBFgQiW60wb/vevQ5BmG9dNFWP4h6MGj+61EJHezzTTUL+nkFu99RsG6aA03h4
7J7rEORq0bsJYbROv609u68Z1Bzv1WZXd3RBibzyVD0pJ/XfvuS13ln1Flwi3rrKwMPD4OxtMXGG
IgPLT3tED9d405c6iyIsObS/aHcznRFcunp3j2QflEf+DPi1onQ6nAb1XO2Rzg2kac+H0h6GAvb1
tLGi4ULyT/GFLQps1PUVgYIa1CFGkdA12c1yseiGw8jb52g7VunFWRqXGXhn8ENeV0jmDGmrj6ao
lyEenpSIJwsUDr41tyWVsNphjQ22tmeuOhbH/XeRRE+2kRsh+l0STNZcxqX6KaEWd1oKeDl+SRzr
59IfQawIMljCJF6bBNcIXcW/1QkSwr74r10AlB8xWe/eV7IJSgX63rHZLa8SosZdOIYHuqC7HGM2
U0S0OlbLtujUDGKkgK+cqBxqMG26w5g+wWWitZWpa+ThJHGcdWB63Tq+1XihHrtz99mQoAo43Xi1
i97zDn9zpYDssXLM86xuEa7pGqzXm6u9zHrTrUIcmCAHPS6ZWzxqnMF3EfuQ9GDxGztHAfU2chKQ
Z9XTzlTRk/1OqnXkMaggoa1J/Laaac802ajtqdvjpS15y8xll4yv9FArMIafVVQ2m4iSwH4cFMC1
vznAnxhhHQgmj11MjlqGmPzxP28kF+cQn7KcP79vHxS5omVLCPJ2344MPa+UopxZgiNvqUuYbjun
NyWl1qs9VG3+M2tKlCvcIaxbV6LkjUEWB+ZCaW7et34frdLcQ2gN9OzQqeLXOdLo5JOTplEs/G2o
Rl7znm+UmrFUqfbJ2yalZFueqdTh31WSahneBzDNw3hRfNU8XEGBFU9S5q/KnbCVXoX2rA5/4QoS
f+XUDXbUfMdJz5q6yIeUlrTtJ0K05842kQ5WT014/E9iA1AntYgosVUq2ABXqB7bf1kCaCQ0drqK
PgTavgJ2FPsdM6oaqAr46sJ13/dOUSV3oC6NhwyHky6YzUkzftiOGS8iXxzTt/5iiITKxiRi+IhS
6hRzwIhTbUdkVfa5oWqwlLsobEusNjmU4LJCabKw4kQMXOP2DvKPbx2y76XxalYf7tOjUh/6L1YR
KZKLD2Cf+OrhoyMClB9LWS2jaB8YnJKpWr7FLmxICRt6Q8smyeFswck1ye1Y+O33/hd9/wdhIYo9
ZBxD7OAl4P9mp/nVczH2H11TEBwvz6qQ+TSYtbGUNxL3c/pyPcJmW+ZoNjW0Fae1aKWJRzCcDN5T
5mNWX8quzZotv73CTe4sOt7yt1bka3bYmV8aGovvkpaEtPlXO0cP7MZ5oxn7Y6ws0LCHth5VSvHi
9wkGKKFkSQ4LGSLMKBSUhmZmv6Z3YU1aQr9LV+ugb6lkM8vtWM7DuRBO026sUGucjTcORWB3gExQ
8M4YrbDzz905Xkzn9A1CsdMAtq0yQpUBtVNZH7l9xKAlmmbvQph4knmv6b4FqppUEz36DbGk8BYe
8iFcVwqsVUDkMB6k8ee3qjLKEZNifbbyLfq0+dEE7rjLazv1hNs4Od/WXp5KRBTmbmHefBJ3BwbH
qFeZV4HtmKm/7r9y1d2jlm2MrCGoSqT8LdAM2DdNF1mnAy2Ly02dU5js97b8+3rrkAD9dpn5avcw
Rf5944cyH8Xvo9eDt+m9JUx2cXRBxkrLcfIbY4nPjaawlWQ3UQRB2HheRZ7Z6WG1XywOCE8Yh0Zh
PpfNiGcBHOCI7TqoVyWtGvGPntpA68QOu1dOd/A7A8jWia6HZ2p5fephBSkf9lxdDoAw+otgB0U+
CxvL7XXeNcoOjwOfQshZpQ5e0z/JaySKzVZxPpZkuTzbtzV9MgDXbSO7TPtMPePWeyumsITqzJVu
VvfSoAVnFi5jmCsDG1reVgyJ/T+Rz1z6Y9z23Ed6ZEAQFXjhPDNJzSo1iKr8FjFT+ipxLu/C4IRT
eaILcyukWef+r4R8ISPu6rtjwgnxYcr0UggVqTIuswHiQlTxj8hoxo4YOSVmx1/ZY7Iean7q1U/i
XzBnsQlqNkr4ER4J6XW9yZCr+lILCH+RMWiNIdXeCjiacvS1zQhVzxhxeYy1rtxHwB75CW35QnWi
3sbJYb1UhHjUVDuHEe/ozD6Sj88yP2DnL0dzDh7fzZQXWErd4qeZP8+WY+ZG+s2HvzcP4XiqGGzJ
+MZMffuxFeYKCHKzfWRRjjKt8AispHpfjVWjka7dGf/i7bmeChRC2/MteicfZ9Tb35pEt8g1wmKR
NZ9jIQRKPINijz4KVbhx91n/ax/unue8BzAyKE+AhnRp4197T9/Vvmnr5B+sDdOyDpiuVsOWUy2u
4SUaFJedVq4xBimzkBFOrUtC0+HVX6dgGgU4WntzIIcd9ab9jpSGRRCh/QU6GuvGS2Y6ZN7PWQHg
gohKln9Xbm1ZtHYqMGwfwg9Q2FBiOGj2hx7+LP1yz4L2N80E/NIwGre+igsjYROnBXzdf7n3xADn
lhLIT2oEss54y1c9x7SdqbH3X+H08Gn3CmlSCc0V5ln6N0ODmlRxsu8waVybVofHuPCpRarr4CV5
ZWUO2J1XdfHttYONBrG+IRdDdiHUJtFC6qZ+IJUw13OGycBTkACiOPyG0R3uMSrvb4Q7QpRBfRZJ
JVUfY+hrr9lQ6NDQqPXt8FvoLDvCGMvpH23BiVRDaoxw8w9EE8dN+Nbk27rd/hcKMHlsg4a2ZSmb
igmAfwoc5Fh6nlCFnnhT2TDiOUeyu0fUpFTd5trnL2r6ZH0BVNTU48JuEyBnZqe4Nibu2S4olrkk
U0N+tpJMJ1nducDnd3/7l3on7XmElN99ojWvde9LUarMBRrpRlErvELqA6n45QFR7/vzH5QjAeCC
EaEA7CXtPz1Kc+tsN8eSUy3TOTTrdCk/GpLzoHAaMzE89LqG/g4HiNJSoVDLoCrOD650yus2v0qS
yWTcdjx/BvOOb71tlcuZbB31uOk+1UFSASlnhnYt54n73y7p6wYF3tz4OqVAlSOmcOaz8DPvCNJc
gcXpbZSQYwcGBXWe4vRqZfi9RB8i0NqS6E5hkocJklnhua5tmPWLeIbOTFrKMrEwF4XygZqwhUT3
ep+87CoILl/kdFcT9phmyWj+emOMbnBod04MZUWPWD+GeMLGVXiB3Z7s4MWx4Y7XGfLHGJe3FCEo
O/riIxZjeqnZWMZ1hP1XeH8c8EbnU2OtQVzpV3qyqTAm75HX+zz63L4hggV1gLyoeCV9XdHc3O0a
pD3s2kPpVs/ckTf+KZ7OTgxgc5qq078csJTAtT5UrDzZdRnZK4lfqTp1nMqKagcv7MrVaa+VCibn
lBkPXc3jkRm97JiVLl9MPuLgNqOivZYaJeHBC3bXfUwFA0FY+0iVsutsmY5+8nLzjx98cSXCnf7d
CmNzUd2a61OWyjwBpfxu2H6qS7gy3hcK3x+4kizwQmdCzprK1YX0WG+yKy4h/G19IIRY1J//+6hW
sqwDjcnq/cQnQ4jw9gpore5yyDaJpmkX+5F/wTutG/eaI6samRW6JxtZSmSajifXQyEiyvaNYK0P
F3RF6363X/5EGScFBJtWaA/2hXbyxBt14NRNP8xcmaz9KXhfCtpgs7UQV9IA1FJDs+lEJjenCe3r
IZ50chsjt5LcIfK+vu9BuC/89XURdCStmCx31MqipGcMmLX3C/tY/XfMy9BajmjNRYurID44X1Kl
iS+Y5RfWpItAbGFJHKZJz3o9vg8ainLbhEV4v1ARfM0gZBx9bl5YIbU7DnHlRa2hCe2SlqK5RQID
JrtIZpboNBZO/lhDFBy0Dzy+J1JZ68AoVvtZuuVmhRVAUPJVMFKAAVEWToVBGd8wiAR2sDxgNOlJ
T4RmZi8ADVDse/aOgV3mnFV8rtkxAVg9mH2uzH1CqEicz9/okqWm3jCnS56k4FGI+bDtrO41WDY3
p3KcDU0jyHvqPbSf4+lAskLehxLY7V87sErgmB93wkjSQquPJ95EdkvIf8xkAo6VBuiz6FOpZ5NZ
ol8q22FadhBiaQ1g9LBZsUkKxTjiI1KWXkAOGRJgxbMP9HTJ8uZAqYCyaNy/JGoC+Toos1Nnjp8/
UG6tzJZD+EmMmT2m/BLCh+5KS7+U6fq8Vwtg7A/N80KzH/z0YIqMPlKHtg0l0+ty/Z5C0kkZ9kHH
FDKDAxE7TmQ7kJX7enGkTqLdOrDP69AyuakOQbPGUAfYP2KwZYpZqR4XDIa32m2qOcxCH6E3vjzO
6ow5lrTE2aCdKP0RnNTCkQcjJ23+zmd770XswaD0Of0mJ0oxZkE1rKGHw06vazVPh6PFsZX+wNcV
XWGdDIy2xkY53kPtC2dbwGHM+CjeH1ITrOzxbOB8i1QJO/Vq8ObRVsAqGJ1oyjnze2JeFrFHuXZB
AtJh1ojb9ncb2J1o7wKXs6jfAYlwflyql+xOeBfMonu/N9RBx9dfcBrIzjAhopBPpfCTDUK+bS4C
T00/1c/s6lwKi7rqVL5CQJfzrWgdiKewSxvmpDttFDA48HjCbLR0YMCvwz5RecyCvvVFox2iioK2
iQCSiR8XqzbTDL4yOAx0FoS1dYRywvfKTU1ibNX+R3YgJGEpNEdspRGM58nDkZ8SNDLz/4iF2Hig
ofVMKmmMjTnxpqkCYE2n75mnjla6PSblJgzatJMhMPVKKPkgCe5zMaGJZzrdbI6eS0cQjFji+DID
6P5J8oxM58DkZYFctbECkIgym0lt/Hpol92FKg2N0oC6SaLa7hgFOrQp0sM/9PJjieV5jgXeWEKM
3rKAZDhRDqV4xIGZ+rS39zWkKsAYyOB26mfQMD97ZEnTNs4U1HLswb+vnLsItgmrp+cuqxhIslMy
TcWV1LKY+BrEsJrooohD8Q44ZFXLPyO7p+LIbz1FVkiFWfDv0yOm43lckyo5ioqjNqz+ssbmWXbP
sF/Y7a/Ui2wa3+ZtxBBsMQmNP3Fd83tbJRa/CdlpXgVVuawspVG3lvSMwHJVEx1Ka7vLotngDir4
UCOGCGgbn6l8DCEjb/hL7XwMsijgls9O6yZPA732s3OUGSSm2s2331NKLWtXY5K4nR+PHm4PP5Gy
7Mn4thnFVA3i9fnfsQyCaL41+LwOt9pzqGWo35YyW4fp0MvsLWmbrhN7i+HtkSpeAl0cM8RxtF9i
fdvxNiSuerBTRdkeCn/GFT9++R35vBjP7Zt7ZztPRIpVM3HzuOh044eJ3SLEfsqcu3hSlJNF0cRv
8wxJPxrCL0b2wgrIrsvMBEHJwcaDO5UxaMBkarjmK3hOnvTEVopYYRIakFKUXR4DAuRSQD43nNvx
EcznbXe1/la6KtEyDvpMC6qX1sR0mPCvSFnIoOzsPX2V6rIbtz0S1oeh4X0OTf0ozIsyO8cDrbz4
cnSRrhC0lozR/JC4JMLOK7JTU8j/tiu7nx5gbKq1TqOBm3eRIQxyFj5P0inhIgIoja+QQLjzfXB8
C2HyQiEc1DSUsgS738efunk7WTsp6cPybgFeTWDy5xAvp/kihpWjkoqtjPD5nkMnf2Dfobaw6KOX
oSfyHcL0G0T8LUT3uPQyyNDe+HzdUsrcEpotRnzuYOA+5sw6nINLGRqWXtTEIU/jBww/qjuQGgqe
0UxZ83XrHl3XVoFoFf+nk8pLl4Y/pd9EEnUkdXvqJhFKVzhb2grvL69PAbEi/m+dP8VDX5MSwZkB
T7ofrqWUZA7vM+gZpQWv7hxAcYI1IuJBzPMw2RRVviC1T3lu5wUXzE46jc01QRFjwqQz6pYQFLq8
9oXSuCuSRddQwZvKH7kO5d7+/D+3qkkm0B2dfydVZU8mo2aqDOKnK+fOmfjMHb2C93B3M3pfLDWf
LhzSj5oprWsvbjD5//gSv5WF5nGutWg8kIDYg6JzHd6rohHidrF/WTeKZ0+QR8iCLo07VPvw3CoQ
XgKV1MMSg0QPuoqaoaGmuUpO33xuzgpx9dgnzTDqRH7ab1kJOylyhCGMkqpkHQ8JpE+rbb4iC46F
Jct3ehBMMzz4kIEFRFyi3wr06u87oOjWsBG9dSsYh7bKu+0PnBB+bLLY72yA8DQqwm2xiarEyaaD
oBTHVMR9JexrapDhJQ5mgpVI4pVzl/wW9CXUDZox/OeSE4bNRGpBCHiqLi2aupLgKp5LRmqpvXbN
mhzVtI9vpoaTSznFEJKro1kPsL8r+RuU2gBkp1Lma4qDAr6VM4AFiQtpcbyOgJ/vrpefn2/Qruag
NJzhkZ5r1gseBT20Wud6ELR/xxKqvMPZcCNHUk2APrs29JcVQmYFye6OvRByKPG/5HJTj6NRQNhp
Y1qaiQ72QLS/7Kh+oCJmFGShNE+BkAElKVJy2kQHkXHt9DRNrcWDENfd6jD8J/CNYODnuWYFM4Xh
TWr//Q92m+fhNF+pUOJGnyrZGwB1XU0CatlJ6/o9vsWZilAyOUVjKGnYtkxdt5Ep/ua2bIrxVQAJ
UoRWlCsMQaRPy9QHjOfsozNYIys31CAsANw2q6S/5Xo5RJa2fmeKlQh18VZYSXhpEVPyk+oETgp9
7BMkDUR4GDCqNrvbywZMDMJx2WavAsIBwEQJrn7aqVMkIvGo0zPFRrEldPCbN/a5b1wmAb897ZJV
mv+0AKXcfAYAjfXtPvmPtJAIkWjU9MRgsagmnFM87jSgrAxKtGcgCbYMH+U1UdIEZC0RvkAC9DUS
ZWxXqAkDH9vPHdFFRo9t3Wck5h0aVBBxkDeU5pCoCgqaEt124rk/KYcPrcpcNyBr003TWGzrv/en
gtqQeTIYWrxT3SjkmPdAPjwEU8V/dJrpK6SNMvXJWvknGx3MYDpT/b9ekgWGc1g+81mG0N0ylvB3
dJQ84Cuo8eMxMGIv72sTodh6bbUSttzG5WuZcyywYvSxurX/M6gUihcmvU+OM8lYl1njKqpOwSwF
hP1aCA+Hz8WGgwD4P1SLjnBCK9usykTLBhclxh5w5WsUIB/1U6M6yApjAOdofn/SvZQe7tyzScd5
EKWQxQM95Fh/99WMp+HreODNzsiU4z65JtcPDCbibG1NeSf4ucOSfKu5UvvpHv2zMccwEEA7AX7b
huYc+e6lvGiIA0DMposR5a95uDPQ64NazDPUv9snZDavNtBcFJpAHxTzRcA6rkxYAlMEYA/0MYZW
EvXrKbf4NqlTz4x+bgUzJucD/7DQ65qWNNMk4TuGSleLfACjvVqfyi3a/dbfF8gWuolRTmr9cUPD
tthw+7o69U2QqDD8MUPBm7D3VcmdaTnt6xiWhGMUStaC314p1fmdzBJYR1MUOwwRRZkQj1440qJW
05L4YvcLRUxs4IDGHeD/nxB+F+rSFVBRqjPNd/o36r5aUsDB9DT38FUyozFBaMzS0rglo1INqVON
JNWrcQt1JmXs5aysX3k9SABVaQaEzJY3s/IGdWPL8EvpVoZdpk8h+JMZ3tma2KzPwFCDyVZ89DFJ
86ctD96cZSY9JghA0qRB9IhJqrGEQ101D0GThS9FvvpHIOUG1BxQj1/SJE0NZ0VKuhFIFBJsKUOa
YG5yH5CfFnl4d+nCLnmSG+zMxEv1azZcmi0vHQrkDfGtXSgxDWCGRrXOUCO+e4/rTRBbnhIpQgq/
eoD1NHcZER9a4ukmART7bSDh38vh36IYnjzMkExGPs7L4aKVD9GswkAV7+uD00QTiU8+80NP7ANX
R3b73GYIVIb36IXDBtTzm/ebkGP2qL24D6dksNn8AiIMipBxWX+ooiX5gQenwR/TM4LK1ymqBpru
sfMgvg==
`protect end_protected
