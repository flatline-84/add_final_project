// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:06 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hnqCtILs1JBR3p3YBrYNreZO1YOCz9VDXnAErLaa5JWhJcdc8Vpgg01j7uGWd9bD
zYpVvEJSYQsPC/fhoFLen4Boc5f1jDkNN05o1t9M8XNoy/PzcreKBKY/xAkEds/5
yCJxrQUl+iaGlwK6wLofLMKuABE8fSjictpE614SvAc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11200)
dNB9Qdw+DefmI98c7nYGedZjevxByjwVxTuFcPEzjSwkY2OvY46cbrZavNVf9JBt
b03XDp6h5DO+ejrGxtLMvRnIVhpE1n86FxPNhEEhp8TEZzyEC5CT1mDmwTC2uCuy
piA2ecBhqsMe3ayuQy7an+9k7F/cbsy2cOwvgY0zst4BhiiQ4jgG3XNG3BpPjIBM
jFK3yWwqhs1BwkyMgOhcxHxggKzadvKXaiMAXJjV+chc9uTApBKhGLKGQcIBgW++
yaetllpdXgZ8iiZq+l6Wo06EobeYYi0Y0w+k74xv1fK0xjN9x0UGAWgxwt/lo74N
0vOc50VqXC5RcXmsya1W8OFrZXf2IJJzLljiQAYTw07tHrjZ19UCTCQrVantWWpL
kW32fl/dmr3X3ZSbOc4Sz9sPvMlaacg261oBBFPhvV8AmEQw4vKeSZa9p1L7wcn8
Ijg8bVWsPJEZB0OgnX2HwMYHVNm+bTmgvXKrneosVtRSEKeuQwCaCDfCAUoiEhng
8NGbfHZa8msduRbbLDok5KXJLqSe1Vc1ceVl+MR1VLKqJvnmrWR3tIbQ5vmssweg
RJy191Eux6kRlzBxB1WNNNSYcTFuTVLUgNLvbtxM4ofQkYEOLWIWlHuRYKDIK+21
j+T2Q/78ZQdc08507bQIo73g1NnhAG1kCxuoJd3D+9iEWD6i5YJsCKPhNaTznRa/
8oW1BTemOdUTQCxfKAXhaJkSQWvu+McrGAGkDM+h0fefTZop2kXFviKxBoj2KJfg
XrTILPlrtdesVtm191FD9ONweqNHoDj3vezDOW6BnyZM9knBeRKsFU3ytV1trj7M
PHqURpDJwiQtei8R/yIiapAvBfGdlGvNpQee5w+kN3AuNoSSQ5auMW01W980/DxI
dw0MSSc2PnOf1k4z54l4zV0xAFpAqF9ju3nWazPBHjtnuGhn7dAxAF9k/TovljLk
awKzq6UfTN3751CTcQx1K1w9jSzQzFDsrAJvLJ33M1splp+R632bPp+H/i5WlugR
Srn7t2svUdc5s+kYnF69XUNPIMf1Agq9+Gfd3CmdiI95sTQAtcjDz1mX7VbLgaj+
80fa7q5dxCeLlf6vgZiXsAl43Y1PkWUnNY5pkvJbk+Bg7RomXD+JoICYpCOD03gI
2a0a0wHtMJT2CuKrL+huBfAjXzR2rd623X956XWOqEgkq9YFEqE3WUp+5IfMK2wP
sOHOO2pCdyZc2i1f5Kgdyo2iKhrrfJyIETYsAPE4IRW1DuawNQsvqr58n4D5wUxP
mBzwVWUggUKEom9BfNEPIw1k9Vs5TetfqLGazL6v8PphOLv+MuueTqNUxMxLFdS7
pzM7FbbsKY2xAShRPlOZCUDt1Fw37l7XWEbS1uE0gH0U+Yg3XXRNbeEwJf/N3ipm
ZEjNSheVI7XX6vYD/apwN4gR0oGXpUKi3FJxZoGB6YhmdoWtMkNfWrrfMlgMc1q2
z2z6ZNfzUJBzZjV0EqY2tcAEb4NHJ8E1jlhKHWe+vU+QV2daun1QjHckejy2ySo0
4q7XaMTfFqy4nfaNt6XpFwUoZRmWL+J2MUAWU/BNSr3DAAu+0cUVLtN0g5sno9PJ
+Bp708TECBy87kaqHUm6diUHTlGxM7+4jGprOdi3/xmUFeMI+P+JZikYyxm0L6ng
h9vwlgYc5F+j7Fs0vglPkIH33/ato1pgIJo1w2YjiOfmh9ovZ5tGwGtDdXu6PGhW
L5KyBiCKggEVuQRP5OUDpDmmdzqVmCBVC68QhdgnpdtVLbjvDRdkCnU+c7Kn8vQc
Xp020g3yiKQdXJ6RpZUOhtK4kZjDjKCvdX66E3GB5lStw/HnpB/oDiEu3ehGqb8t
dM7X+5+55pa11k6uSgx3J1HqEjcv+BhGNtQ0tWdJCM3qtDbZRLhE2ncPPO4aIfmD
+QPHB3t++pLBvccEKKYjSeBEMQrn7vi8E42zhE+xOrIhRjZiNKkj0mb9m8jLoVeC
GSqZR04BWCunWBPo5/0vTeRI1eMzw+B+7c4bIuOKyO9F94Del6Y/DofKNOxBkPkr
Fot1xWM03OdHnwsldMsBq64yKSyA2PrMc4wwB5hgohuwgtQJ+KkNhqqTR6uea2fs
YfV9Ox2JtAMNjFFwI2X6wxm2jAz47dqxfrtA9Ts7Ph40t9gZGMr18Cj7eakXOIJq
81e4XRXbxclHJx5ScrX+Bf9SpohVTyw/Dc1kSVV2KnYetCOoeiLzsm6vvu87WDlF
WYRQjBxqqYMT6idrWENZUbAUwso06XTstazp0Wt8bdi7fvC49OzZK5SlXJBV1oAF
7znQ3W7V5djpJhtfBiznL7uc8r2sdICHPOZRWo4652ttIAt5dadVYgavAhDwg8Ji
bguUOuFxJS3HxV5cpo/20kkK15iymsTJhjWXUHksw7RgTE+inGZuZsG8eNG8OZKG
6SWSF+jeruad+JS9mgV3GD12G5rUzDxfNY6CSJc90m7gwAMGlTgY4G2vJAs2kO2D
63LVj08B2NvvygaUjbq/rYnJdaWM+YV8n3iVNUd22bZyptMNZLIyl0wVIty6GVZq
nmuOyHJNx7TX4i9OJ1jcx7UwFSxDAcpZTi0Y4aWeDqmVVIG79rW39A632C+HlPO+
FEgDfF6ml9HWT/Sr+eipeEfb708jn1ABRSKikUqbb2D/QXDAchTcBLMZP7uMOkJf
JjEhhtItnLshuF//uqY9zUUJkBbCnjOqMvTc84yEfr1pkHGnC+wj/ib0hG+M3XhX
UJtUR/E9AD22fYURafB1CVjhMny3C0UCe3mPHTENAs/GfpxzaFHlEGGBdM5Z/ikP
htCw0RvzJKTH/KfEKddcIXLthqaUOE+G/m8Yn8rqyXGEYlSuuoe0b6OIKR0Iy2Dx
Bj1ICMgPyD3biOVyMVYsM3jhO1JscNtYtg8bjRupRSHCjhJb1TG8KYZBQQeSuyR4
xZzMfbEfr8W45VQYLkKh+NACtXQWYSMAb0CsNObsoj6SnnHlGhUl/aN3O4t1kUtn
OltUTgkfP9iwZIJGMBN/JyNbPcUl/susOkn5QpFaDPKRcKb6waAUFf3m9LCf/9JG
lJ6R15cU9NsY+a/UrLPJ+t3aaeNtFlQnZxBsOIo1PNiccusNgcyDO95/pr2CDli2
OI56ce5CbynjkkZkhXn2Myn5s6lotryFhZ+mehJ2Zf7JrApLFQwkPfE/Yc3ciuKd
BVa+Lg3zbY5AHoEDq8Xl+IgP10Cp6L49tlUr0KvNDMFbf1vh/wWP8FGsI9xzZSCo
/zKPQ1i8RUZ0pMsHTaDfLPdvtoTNT2suop3gzFmlyd8C5iQjB5v3Ec6rb9NhyZIq
fBssHwveWcqp3SuLeXwn9QM2EeVqxQ6A0IR4Kx6R37wNnFbrfQ8zz2bbE13LDpAB
pOdK41Oam0pWButpEO7MN2l+GOVX6vtmWP8uuBw30edsHuULAjq5lJl1b0mggeLF
1AV583DAO2N4chiAAqBDcqEzBwYmS3r9R5WQ+hQmJwkQ5gt94J7hfVskiqTsgkwR
gx1vmpzVm20OqJlKHiTpcjSGL/xXMULtsDGfBn3HMJc0BVWZkZmUu4aRZ82kyk3q
lMwLuZwxJwsDmefXys2dsx6MvhmyjzhAxmBP9h4e9GjM7dlGcvAnXVlWJOmDuS15
2FZc2lg9LT7UFN2uhxllB1hjXDluHeJYVxxG5GDKQhhLpoq0obpYtcCh0D6gh4un
day71Nr9BK3mlID1z+4vY8UQZJ8laYvLtz8Zbh6X8Y8awdgmCkH5iDp4QePSYxwB
QzUQWX8fNfFGouwIl3x/7SQcf0YVdcAldVMAOebr+/Jh3ufeaSWFpsqspYCvdMrK
ND4g84yMQTnkBhzU13KCtP8OLvf/WjaYrfui5fWi4mw3Fym3Ln/d+FBHazdf7pmY
zutbC1fljcmWx4TVdbQNPYIHWUiH8HWQbcOluWLiCqGUTy0IXafYDr2DGmBjfETB
2kaT+zR3DUp+uWciXVKFD10XVW4xFWNg/Ncd+MC+ZquLsGgxwu8IX+JCpsxyz3PR
/Oat1FNB00gGa07bCP1NlXosztN1xzWYcGdaTsC7qIkulDlLF4hDkJoVQxaD1TuG
6JGtC2nfZCKXgR3rv3QMcHuaRQlra7CP7lUwrC31Ddc/xJPiEX3ymltEENl84y6V
r96eyolnbcvBMjvADqGluXD9ttDGWkGGJSyYgc2hy0826A8NlR8Bb0dBwaOz1qJf
IFc5Zyxv5yyx7yBtt/hlfgfoAK7fxS5Z2WIy1iAr9/Di4JSEYt4zdjmBqY2IUL9d
pEAdZQqkanvkuHGh+s0ZRQeIP4cD4nzgzgQu6HHdh+vdYOHdKlKVfb8STYEcbl5p
N4Bsk7ttH7rpELlAV/uegNtOAqH5yjSg3tt/nEE55al/HvqH2380lu6GxU+zGiT5
qSurDvJpo6uHC3BAdnAalbyfQ5aS8ETf3lKkwVmBCNrr5Yp9lUbW+hzfJgNq1Khs
DRugkFenQAXZtLGO01eyg8cB7RhzW56xHhVp2xHZEG6CTAgHwcgAK94vpYt/bVLo
K4HEG6Z462krmaE8yhqCUL3tVOM53/s7h8sEWxHV+5pytthJyGQZnRvY3J+CYACf
yNGL2kxgv5alJgrpchowBHuG3FAwIrgcwk3mBit/wU21XRRzMvPoIk5/iLNz6Gz0
NBsD8lDV9r2zSsYvyskk+iyXwvlnLh5wSH/kh2lR4vPJY07j7s32ox463osTclZw
SF5bXd+wZOjfFhAXeIpXV8wKoNKIEGDZNRNpMlN7fhx6EnVH/yIqlr388XETv50C
I+PukdwY2tGCfazXxX1vkBF34uvPG4avIN0ftipMpMk2WdHV+vrYe+C1CaDPQSvJ
rAiJ4UDhSSSYRuQX3aIKahQv3+SIJyyYfkoHE7FAB7IvjqJ/HrhrTeRQdIvs1qj9
Pe35/l/X2RcJdIFkyyEYww7af4rzCOVg/k81kRg02R/nGT7cDv2wYgDW7pVZKNJF
BC+JWSPUSDWElCoRV7atKlTAuX1ZfcaTa1NigCm0m9itz0nBciba00XLARhsuPjG
LPiVwBvIrRLsK04EMlLnevEff8yA1y1ZzTVbZQp53p4B+RRVe/993rWANmGGg29s
DMQOvolWHAMFSPze0dVVu6wHJRusNJqaInzOm+8I9Q9cwl9tvybv2KaLq+pUuTP3
7iXx1KmeRUggMXbLU+8WpO1rSRLyeZRDFc3eGx9SHtSTIKDccXp+8LDsFjE3glWk
eeDMT0oSv4awwsQi68sPbzQzLNf9wuBUUCuGL0VcnRMWBtQ0IzfmHkfS4PR2lNeo
h15pGN0dHZmI9MnPPF1509qohWjkiBbEj0SupII1s2AwaXjrqm11r+p0QKIQidCz
aLWxJMB5LJbHvBos+bJ2lB16xwyYcP5DCvRPX72lo0Jbdn9L+p4xU2ul4H0YFZa4
p8lvrVssyai7sZnWcPJDjqH25f3e9eUFTAfAfn0rxtdJweGloU/xknv50QjfyB5m
CKR2odxtwoKwW91Rddd88MBdwO6J/3Ub5tU7fU+MpewbFp+3qulJnWH+CBVlMpj+
YoEdsIhF6X1H/eWqO5v+q1PIgv3bU9DmMvlZzv8QltwkhXZgKxSzFcNYKd+kTPQ+
2CF2aSCypx78zgZ3QVy6t2WiU1VcpvlM5aiGZsIncA/RpOUMyRtQV5at4OFBWT/v
2mgR/v7eaGJhtyA59W1IlZBdOOLaBwuHy4YA4dUnUEu0JLPR35JXxJYgMxPzcy3k
EeceHcbqBWa9vtuQJS3SXMkNtndyMjLdDOHnyxWtVFNUght5r8fvKZvq3+IKpFjX
2ipq890FjJHv1taDRpZuP89WA9yMBywWoR2eGaCJ1BNlVLTmgSJtJ45PNl4fMTOM
M8wyFbJQc0c7PCDZW2pc8901wQVmpyaEjTbmzKKyCvXBSc6QpLZS+fwOnNYw/xzu
abjnV1RmZKOHQy0ysbPbHrTql48BZeEtMF+5CpwEQdHxed5ajlqrCKHCyuThxaL2
hrw1CS24oFE/n/o6DJyAyK8iFxbpGIKOVCYkRIYDQU8UAwsns1uLd57vKlCIzs++
G9UrwoFu5T3c29qE7eZSX/WV74o7sDDewQkAUcPbwJcCqfymy7INC6Kmq+yXnUX4
JO4iTHFeTdUdvOYkxA/wrOoWyW2I6E3QLp86SCwckBBYO2FZRvxc4DehTwsXWIXI
j3ZQR0hR8lkQtXjcMFK07NMIR+OXclBdOJY4LufuGm7a4dOsckQdtPWFigPtA8Gf
ICYvPgZ0Pex8uVJhFwB8xn1+S8sQPeKWkKEMqQLfMftYB2VRQJ970VCiRCsZBIr6
BChs+QhSE0VFFkTuhikv+LLHajwJhSP2kbNIJrc18GI3LfkH5JIOKpZaIccqFKm2
lo9kNqKqtg1uFMw59vks3A6ab66hAj9fon9gPgUbRI4h7xSWCm21OGle6XvfcrIP
AmSQQIhbidwoiWEHrlnAOsTZYKp6pP6FFRkSGL90EFkv26mgRvAB5r53mfyvgIE7
Mei6xTxu++f72idG4Lbvf4lHtruE+dBNbBWdUExATJcx0McsVs1yPA9wUATEIxQ5
+v27OKJqWqgH91Wjg3iRvSQgrkWCBOhhQHXzmaqFRZe6tQqUL4zQXPFeQB2rtUDN
XoL1izTbqzvD7ZRXZw1XgiBz0t23aIB2BfAtcD5hGC4PVmZTy92JAnZLuFR2VnR9
IBLrXg13qsVrOIbin3MZnAKqwERQKG56PkPOfjtWzttVjivoxY3EWtozs2U91bwi
USPXrOHMrY6JtI9f/WaNkqIuTfPrM+kGUav8+Owu/DYfXOjP95gtQe5/r0WREprg
t3KHbGYU3/Cn7Q/YN/jFrGnbyc4HBpJBHc8mzTEguCnsLMVi07ShYfBe9RrtVOaY
VKw0dbjrmmBrG+8da9WAtBplFIsFeYhoTFW5pZCpk9mPn0claJgH9yeXcEE4jSJ5
YAZzWSbPVc3ez7KCl2s/OsoDa3qpzHUVMWatI7SgaAiuyQZ3DJKH/2a56AddfqNI
iZMdWthD1u9q6vmKyM3/HhHZhDflCk9t5WiaLSksDGAW+G1MMi4HIwcPPqkN88y9
gtFUvdCTk5Hs0XxxsziUJ2lf/Z2qhM/ggoyYKQA4a/wRsnuWs/VUY/qo8oYwGc3E
Kn/iVPdqG/GQK7HnQzbT55U9o6VBB3UJi8xH36vcLxkUomJ3lctKm77CvLSYHgOW
N+NURSGhq0MGcAxGIjyHNLKUlv+p1jMDj6sPM2P8X/ZIcGnudniOMJM8nTD4YDAI
g+qTtC3gSI/0ZBVKLFcSyBV/uE383S8xkK6T1Ih8kK6CLvr7iW65716M8OTasBPm
PGZMqOOCeBaiIvE1A+pTxhGmM8SvmNBYLDFgkQzAr6FJYS2QcXEQ7uvaWJdvopxF
6QRvXst8qiVI1lvPBxX0J2odHH1V6026q2BdA8294Loyk/R8xJet/uVWB7wZ/OwM
tJk97mssfPMeAXk+DmSH1BOQXWbao51kSsT7z9W3FGBr8ZYX5v1Q6Y8LJz5DOtzR
V7Z5xYhuakOkG3JoQYXo1wbXgu0UQVfSzPZALX6XyxmAaLWVr0v3AnJLUKekKJHG
cpIBGGd/UPJyDoqC4rHd65/M4Oyb6aD9xOsEB/mqkocpOyrkTM5Dn08WS8jFOTt3
GD7OwMH0n/2Hyz9rhNbIDl27w75y37LJ2E1mkS6CR/wg4NCzcmFwhpsB0GwrJ1f9
wBQxt0XX80gG5L8BoRKVOjlr6MzcYRDwQEVAw+55tEkIWeGSXw7yYPmh8vLoLiDZ
7cfE2Y3PVtEXyv5nVGt244VQsaPXnGHcqoXDz+bA+VlI8XVhotU5PPb8lFPAPLdw
ibPSfVRw847m1sIB+h40oKDX3LuwvKE6vtoKF0ucAeTi8W2GdYrEwjUv4WJdPubv
QcGbnDV8cfH7qzL2Dfo70ww00303+4hOmpHuwOWLhSosgoax8aM5/Uanuvc16rMl
VyykciR+tDYGTwBITCj5FUE+o7DzKeIiKvgMDjqLTtZR9qU1BAb/bpLHRIVaQiw5
LgXRmSRAbQHy9xvYsda/Bf2AALMIUH7WH4LgDxB64zjzbm6MRfqH0/GVm0FyI9Aq
vclKRSRT6gNcgwYtaQ+kSv4wN366zxsfqc5D1FHsxOhcxhBXrC2MYm5h/VjcT5pS
/Ax4DhIzMb5g43KQ87TTqtp4GHWNKlvSol/njsTNhXJCjrOKbubOU2tu/+dzJii2
ndOu3SlER8c3xuLrHpG/bMJ6i9CarXfEBIFIRoXA+Vvkr5aZXwhMVNen/t3Q4jC4
WXE6Ma9DS01olbDBQgklR2tusrIng2oOISFIQx3FcP1xugPkwn4N5REvk5/OivxW
ie+sTvrEHE4UrbW6kFCYLDlXf3YpRRWQr9A5WiAukiI0TP1h7gEZxrAjZUf/yInn
GJapfD+NZ/IxaMtfBWWphxbQ9sSIe4SxEHDpp8x/SYRFnSMnXcH7GzLWb20HfwcP
B2uhdPtAl/KWjm/6wy2Zj+42Xm7yKvMy1iKMjFZ8JrUn89BJBFWGrlPIB8TPZU3E
O4SUM94M06eIABfp2nQOrszKPNgv/0GteXR8gK3mOZthA2hM/BErdC/j47JnMgXg
WZpjma2Ii2Q3xNzWyjVfbqHn1WLEYq5tJcvf2WIBMqcfOthfQTpQB9Q3KpPicqzo
9SCX0aLIWoRXJfk/fPraWiZ4GISm/zYd9OlYEGglqkk36Ib3sUrYsjbdcXs5RhsG
CptBPlvj79VDKLe3uyVOmidvFSoiD8KFqw2TODzcLFvqpnJ2Bs7y1fubMLCNOE+c
AtWH8yzmLwQMDo8ipide5+S0JtECii6tGWQAHE1fh3BFdw3aUiPxnTXi/i2DUlHd
sdyZqdU7dL/CGlr0rKaN58Uk895PEHMU50xC3hiUhL8MtzF8FK77K7iCtPbNBU5e
DJDcjZOHHFTeU3ceQlO6NUnKw8stZFQgJVtIDo1QyRGUt7zWtBz9tI8eUxT1b3AO
xfI+GEDrdvUDXbZTxB/I3b7DofSdojA1/hfOL7oKZVe4EcFKi59TKIXviJA71Ln7
BDnLL1qZiQAvoHq3QGrp0Zw2C0zq8ACYQ3Z1Vpk+jejGpw5srkZGG5SgvuEl9fdK
15LBOEIvvzaTyS3/nid7A3CW/J3k6T7IFltEG1cMFjoyVh9wzgUyZyUEnROpW+Yh
ao5+I0ZIhdArbsXRZ3+zcLsgLl5DH7kaDENXRkTo5MqLDfmpUPfCSomWW/a9i5oa
eVwFoO1SAhYaKwDX4nfR/FSAp5AlezZvUz4mcJz8XDDvrzGX4SFwT4eLImI0OOxO
D1GR0jE/0XIVfk27e8zeEHdiLTQB1igzO4WVrtPXcJ39mX+vzNHXi/rQXDzwJNTP
vnoSAfJT2THm1Klt7ve5j2Evp51tp4FxVrS3GUi+cKSXajtL3EfrQJW+5UZsvANy
/9o/omLeIGKoKZF7eBVoUcvPcd1VDjXn12e+KHzsmEVo7n4XuHcAAFLktEFl8Ifp
PO84A6KmyahXT9SfZK9cK4Pt9cn0as3TS0XUa+iyMsivemVBwRhcFntNmEKyPS8Y
xPT03082EXTgRnV9/MPCHft/ukFH/ka9fjsZqx3My0E6w2TSggN1fPehMLC7QCLn
4y55pVDuSi/GNhSiAa1AkQQi0R3q/H0h8Tr4hNlK/lLyAJI210lR3Ac9dNY8dN7N
kIEHIcLBxcNYmezxUp5+3SoicQkiwLmYJ7m9+cCiXc9rAUcohPqAJKJjFN2uN87B
gyDvVZUnBuWSvPpzaC0PeqI1rMwwlS9BqJaI0RrGmqyVLXSLHjzqIlwVeW5ToSBx
cvaM1kYUycn9ARbJgZdfqu07PnVJiO9CwtFbfAIAD3hb6hs6zvcG33xsCfZDRCh4
IzAXz2PUGrkxI4KxGKEsuH6LxlDbxJ40KebuwcDec6lZa4OcSO2xOMtDH65hWQ1P
SrljYiBQ09qlLRhg7VrtHX9Cx7aLIqw4jBt3OKdqsYfKEMtZ8aL3RwAwUP//5v7U
SssnosEEdNJD532pFvdC8eE2qW4z43E4d4xtvJa+bxjGp3I+PE2rBvS5YcQ382RJ
dD3ultcFJIT+CG4NS9IU38u12iTf7dcVj5MFt5wVJm6TJKXtA1NPoaGuH8oYj/TR
fCG15pnLBnc3vKGVzQBRQj/h7mASro+L6s9W7uWTgkSPAo3wDrtOr7dEWaPG2JKu
q4IJk5elQYUqhjJL5LMzErcQpfpmVQ74wZ0JlJJ3NlQ73vN0mz3Wn7kwUo5mj0HO
K72khpnJwFrm+TyxaH5h1NoCHC7bZtjnlkU/4BepUjrh2M6Qk2NtkQXfe0oHD8Od
e8FwpmlFzL3UI+X7YH8m8e2GaFBySu3lnSiOW/Yyyk/DLVDYRsNnoWOAJlh+Nz5o
Fhs7qpZ5Yhcw/xnNfo9+JGJuOzzWnjnNqTKFIZzaJvvvbh3hRUq5dsJRLbD0eKdr
KKU2f8F8H+YwJFf0XZLDRMV8OKvz7Bacq9XhGkM9AKaE06YTwr4A0jwC4RWIPuru
sU9EFcY3yR4RMvK+BoTNla8KrVo1PsuZTRPJ5A6Z7M28D1T8KHPRrIM3tSopYqo7
ZZh34J6fdHoNWL0lgzqPWtEhQ8GcwwSDM4Ja0WD8cAAnpn5pYjkH6iSE5xpUExyC
vupUGH32UL9k+cfovvdhLc9gHKLuRusJbps6toE8uQwlKdY6zO/EPHCD+ZKuMyls
o66l4MU+HXR1xLJd5Ie/bVNavpOKAUBUdAQ5G19YzgKTUuOHJWpgEVYT4FcJXP18
TgBqUt59GHlgUPUI6mFQzslLvvLfSyuufnjWEmKpQsEnh9i20NHCJF6yEN7o6lwl
Z6QjnywOkUOdpWZWx0nTErioXOEnMdaE5K/4N1KzYZoLKKJefJ1nOLNCK/BKS5a+
Z5aD2tPJABiU90J04taa+Kgks4Mn1TLkeg1AVk1tcpKzTGsB4/E7EciBF/KJdYfn
jP8K10nHOj6AqdOwYwJb5aKSt+8i5YZbsXMGjjNZ73K2kCGcFMlTPq1u4EKLkPpr
t9VGtvO1UKGlXsskzEbftiU7AsWOSjPzS9b32HSulQNhU0Vd3hBFDB63HXCke00a
gWUprQH9qR26kOKGcWkuqz+4drueHBsbRRSn9iHvMolyoeDeHtxRzxlcK8TBHqYn
uBkwdps+XVRV7zGUNEl4Sqj7VwU/usMOqijZXApCaOiZvChWTm0JfPG9scSiWTmQ
568X4+7YiSBNZVbFahHUUHZAUf4EaWTzXlTnyqgh07oyTSRqNSzukY+A4X7D8d41
ME+5Y0NN3JoLYs1hYdnBvZzK+u+ZFISaADhzgCY0zWKVFv1gDPHEDkpM/Ug4v5P6
Qw2z02tald/CVNr7hrbmyXD8C41giXfxu90rzVCb8ce6jSnnRosscx+luwPW2mq+
nL0HRFU0lJvNjG4nobSoaelm9YuL21xPkTuph12W0ImtgNI6cT4S3sV6nEoF03Vv
2vBETNorQkhDfoFYZyKM1SvG3TjYkIWKtp17EBmqIvLgstkAh8ckAhAuyYCypc9n
/RY3vvONkSyMrytudqbn5u0Lxju6Dbmvy+6Tl46JzKrtJRAfUw5NYe3pSovtxGNN
TM+IN2l/sJM80+PyVf8PucRTh5Ho5SOMdSEiRvZ/vleVMMH16GlzPoprvCfEf0ZP
WIrZSIcCH56LoLMxszJ3JsfVuZw+W5K9SVfgaSW3Mi2tL2jVOgpXJd1HG50DvYgR
jZWJDJI7jl2afAm/R3WQcs5sxxM5+9evimfxN+IH4oyZYtlc0AnmW9rUasOMhW/p
hPqZSMx11lV8YRr4S0YqG8yVfTv5qLR96drgM0tyB1qvf1/CYvt4t4DS+98Q21ib
az5YlOFQ97EaJzmp9krEBYqFzvXcO6dx97ewWtRI5f0EKzEo6xgqZ6JqrBviLDT0
vGwMb9p6Np6zD8n1ODP3VdY9LwITL6gDk84ribIElI0is3+93La0PM/vz+E2wQzt
b40VY/WoD/8ZZ3U6svDjwZRG7usDA6TbjBk0whFOJYw9bwJrA4rT9704Cz4cGZAx
xBnj/qzSw4G/JYmNRHrBV7SP9bS1uRIdnto+ggE8t5nLf2FOaNucIsY9gEe9w80m
VCLZwu7YURBOru1QGqZGcLULFwwCZMAMeP2cQlQqAyfPPy79S0fmMNx16HGqyXdc
qSRCgoSR6jTcTNNzFTTYnK8KzKDWkd2qcstJDYMbATEV4TK5nAumJzGdSxxjt2EE
1DmUlQrYt3/943vFrbnIFv12ZTvwt3etbK80KF2717PmRSrKiloiUm7PHHDuyhCg
4wcnbQynUQoMdVMOvbmGTzBhq7hSIbTIsEnXbhrrVFB2wjmwpq5hxJ8Xcq/RQ5ye
6m7/ZpiGPKIdbEoMTtDE/aNaVERXRch+O5hLu9sN1Lmx+2FycDvrpQzmhSStf15J
QSVMkvyWzRNFrOJycwvNPqeDndwI98olAfUM1ITaiWq9WFarJZRdroC8u9Y3Vkx+
D/BhNupvVbkVkKnxMLn36jZM26cT8spDlQ9R4GDuya5orcyzGKsxzTZSx7cD46Cl
b3gxoIA8XifAf05GPIakNIssrYHGD3VpLEGiqRkYxA5/b7v0Imrc2u5TqkNygSn9
syUgim40HptTFZ9dpajC0vh10AiSsFSmDQFRStPD2jvJCiKzkV/gJmWa17ojFn9r
Bw6TC6T8Ou/lHqfnlt7HfUN5yhklMa+3oASi3Xn6/qZfrSuo7NDhcqC3jTtBFowL
yDnvoh99oLVQ/6keubfOjyp5J1+ml6oVxwsLIhTk6lsqLm8zkoUsZZXaYtQLjkF9
YOsOr8vfiypvi59tTno3kY2dy45EE4G4IGBGfNIq3lvmRk2g64U66pstqVENz6vz
7iL7v0eGAMMby1ZGHRqkJDYIRY5GNwX9YmrwyiV0yGNVHbCYtb56y/c4bQYp9RGz
Bg0HSEAr243E8SV+ysigPqWEOOpqhmUjOxunKsmWsboFBIF0k3B5d4WAXlSjZQuw
X0LchEN13j4DNddiY920vkUhPNT+pTJf6YoAyM1JssZdrKmLuBi+oIcDIh1SmyLx
macU6Tk0msgIxUiH3fXzlfdtYS5QKAraRob9o2ZsTQxa7jUjdcb+S9D2tMi6Cjs+
UFG8lMkemLrR+W6/y+FccJBwNUsBDljJqj5INYwMKORRUPuQ2nExgjq0vAySfFLy
n/S8mJTCWMFLIvXuUAlyndyoToXU9cSHV6ch+072wZL6ovopzDGP87JqxvvqIr5d
BWOr8a6KT5hYiJAcci+VZX3PjaYpDcpK8+OKz5pd6HIyLfCQeZfbonpVslgSgZdn
VkJLE7kdkm3xeoML+/2GsF2TXKFxImg6u5xKjuzKQG0eGZ29ms68OeOZAd0ysGX1
ZtX0rv+HemAbNijKfxhBprgVQqfuXplXsoUmOkbgU2rsDbHgSAzpLwJP7Kim9KZY
sjpkLnnJ2P1r8LQ1wQ4st49rbREd4Df/6cO0q4KepuIi+eFdxYTEo9Y7fEtaA6RJ
Oi0gcv80xfH88vllw8m/L8wFxn67KHOjUR7CtiyyAEEQOdelOEKpYlJ5EVv7oI/p
3FQAGbfi8zqSgcrFlbK5FNh/IFAv0OHdkk+L3hEj8YtgLGvBksR/ar+CHPHmn0ue
R2SnnKP8zNK5a3VGGSHTbjE3Pn6cjfvJbhaFgsdht1UBKt5BFQM3CN49SFe2v8AG
6QUOC39R00keUeKNPMMirBN1oFaIJaSJbfjfN4PS+AYr9G8I1nAoVf4iBNMRtUtG
Bx0CTTR6NPRXW9//W0ovhm2NBZPOUriaPNw2kUKvVMkGjTq+e8XitHqZU7LmV0Kv
zZ42+Z+CHB8vPdADm08vuhuNYbBS1XDIcE9+n4NnjYccIID28eZ8hDd7rVL7J2xl
vbvtny3GEr6sC0u4q5v71c7VnVPD2BHKAhymyAdrEUzG+EsytZunoYUHAluNVhNY
MCeEVH58we5vGCpMFslTjzHT6Zs7B9On0Bvw6fGytf5lOMDzM6+OTJwFVvlcboFY
zFYVWKAq286iVJoq9+1jVEwtmxtuYT4IzrmiG8UFSdfgAI9sExbc1pdhI0rQTTfJ
OldBTkfqUT2+kHn5HzkIMmJ9absdopbjTumFOPV+XzZc87t8NNRa6+Ppdvv+8fUX
Tqvfw980ob06MTv0wCKt22YjCmuxjj+I9gaxMAaBcPLIkzd38xSfpkEk3Ojc8mmi
F+WC+eh3EZyx7UD9LSYZk+xFToBMaTgBA7R992tFs+o23OJp7TP6JjT6hndJDjv6
aTM+vazQSNxa75q24gJjkRS+kT1NlYQ/9NXUzRaxJUeIWLOsq7+x1E+Ar+ppXvYk
uO0yF6HtL6g+T5dmbk1H48Bvpb/e96p8Z4/oxOedbRBanoTOy5D7cONkh0CvHv70
zT2baXegiRrkNaW4Hgj3LmIvf266QsY5NP8GKvSQTr3sDcCXUSlXMJisDLM4Ms4v
9EqorpDlQbsoFQ8ijz550bsAQEgmIN9GWDnahyEePwp0qJO9MaYxw8BF+a+nMKel
yrxE4FtMiGsGsB6R98+gRZyxMov3W2dwtYojD8z0Lj9IgOSXy7kjChpx6K4nGMD1
LkkdWNRUUD1Mc3lzsLdQL+fSwrYaDfmoXghd8mTen/rl3qzbQkqSlH0OWtnPAt9d
gpeD1Ox2p9ZeU+GqlikYVY8pJ2wxPT9scbgN2tkA4/IJFVsmmrPLVaHhZac/+S0J
w4uVQR3nG3D+feHvqxi98tgPExb/mw9wSEa/nIclW3kIvCxT0cxdwDIHMLA6bB4m
VRHr3a3W1sPkLv9eYwZn9sU6B5xV2Ku7Ey6tasD5QUoUPhTnMKsvmIHRtB/NoYQr
8uBr5W0pYF7E2jQJW3gpDg==
`pragma protect end_protected
