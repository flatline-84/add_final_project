-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bqfFqmHgKma1UpsmUrXL6Tj38edaDz9hkF0Y9bFTrjrug/FBjxEn0aFExK802SEX7Ni3u0gU7/QB
aclf4/bHTJCeONzxtbWV+1alrIR00hJeZotkd7Nd/1DydMizzRKsUyfFnDQVVjjtHc01xI9HKVs/
sTIN13BjyoQr+ENyRa11buu2x3xx5K/PsGBMcJ1dmj+rvgHrI+9C/87pD3auVAx43evhLjMhaX3g
jEueWQdQi5TRQdJ0veZQ+5gIpRR0hrds0BE40lb7piSSxCuT36bYN/Jx36KtBlqTGok6Z3YAMBbO
uRF36BnNwSuxe1Iy5gJAf0bR4vcfgbFIftc9qQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24704)
`protect data_block
m2i6lEOC7YZqOodzXkkDiwY+B7j2uDCO3bvsRJrUqDRmJq8Vy+rgan2fQnW3XrKrN/Tvw3NrpMWB
KJz66PPoRr07z28eUqcg2lFZvJCbAwAsgojKBpEtKfH5gmiOY27R7XwFVCEPWFLoWCdetLGWs0L5
tqMw2Edx+gicm64Noqjscpph7HhpiJdq9b4Ch2aZVCVvDHoCdH5PKsABIahCHPaO7TGCH0QyBaVv
0q1OBhmRgodMeaXLmPchT10UmATbrSTnQfxsF0PB66YyeWbqR35qhcbWd44SxRb7T8WCshor9p6m
nBHq/dz0AKACudFtIBRuL1Y92tj0Px3f0FoMg4IhjGKiHQud0kWoHhcQem7BHTbdpLuoMmhki1AX
bvs+whfxNp7Ygue5umqiT/uZjaCVEgmv9podgUXrgfPlHEB0ZW/e25VON+g0zsTpb7WghsNBqH59
LecNbODCd5L/kvrV8GhZvB09uqHKBzA3FWemX4cQzYQBD71Oej+XUwUKJxsl48B8MEj6RLvD/flO
cVNKCqVCfEobNjmggzjZcgqDxWC4Wpi4bpH3oI/KavAXU7m6qq6BsIZ39R0+lV63jIAp6zZSnmOo
n5G75Qhb0+7On9vF4DjuXzpgsqlAaRmwhaPF7YCBUC260iHi4I8psY0OMgoepXNXJk9ir+x2xEGr
eds/5wL1LV2Vx2dQBzGnwNQFoUmcBNwOiubT24OzSSwPUxW+asuM5YEKupeyRj9RysIamTSpIg2n
Qnm7Fv9Ti8Zxx70qRLZ5HteYKpRFtNZgrGkKMk9VxSxh5uk7HDOwsLAOc8aOQTsSCPnftw29i4qa
F0WaTNG0zcatD+mbOya6ohRm6UZKqEwIp52T+m3l6wdX8F9YeGLa5+2geybAmAA0zmLa806IWil5
aD2Uun5lt7HldO/aWV4Gx9Giz3elhrc10JGpfFpjGdKJeQNxl9hQqmd5FRwfswvXIiREf4k4cAXc
OeeAHYBAFNPT9/BGP8fpdqVsWvy89za+yf9wlSlEsyYNWsNfRCbE7nCuHlIvpD+AM8HU0ZhvW3H4
Yluk2Qaz8IociaENXmlokH6kmLfgmqcURiYZIkOBV6nJi8mxOpGA2lQPV8NCsm2iU16SGsolS71E
schViu6HyJsGTIYV2GGkH2nU6zCmjVByWHEY0tvXjpAzo7sHYfT0MypU/CpbEhaMmBl2Q3uS6kXW
qCwCp7teeu3McnWJkEXTdKIqegyfpq/6KGFAd4uxBobhh4sjHaACOOs3GKR//S9W5EAgIDPDndlm
VUiUGBZnPSnWtgsNMHHMoZAKEQN8nM/xN4W5Kw7k31+zHKVV/S2E/6RZxFoZ8t/hOJwPZB/dUmo9
qNXGWs9+cA6irOPtXu9xU5pTHrRqLTkpkkD+hlUP0m0ScEiHm/2d+Zrrew3R87Qcfgr9AdpFoIfp
TWGv/wUsSyz3Qa9QYI6+Ape6U0QV3pxGk4tXW1VuiAx8fUGhQogDIhVb43rjlipGAJ5Q3wN0OEtl
X1gZ2tp/ZNqKkNt7qOPBxjU2dx5426TzyPLBxaVEzK5FC6qJkXibVxp06LA17fBZeXqFKK/GwPC/
j5yKPKSK/FE3DdRx5wEKSIlU6xxjZThOuyvAHsE/GcsJPlIY/AvfctGTVoTpez7kix6RFW6pc5pz
IKnpoDbbcf0JfAP35XpmN9q5gpqdBHVZ2+vlRxyDjnnu9qFSiq8Awq987BauamkGNVfT5Ve2tD2c
ZcZtBMVhZWSXM0uBSCFOxqENVgB2T/fyxKtUOEIxPxXvkN7JdLvSOnklP1UOr8cfYYiduzFkxW0T
+lHSmWmYDs0OqEijfo0FPNvjGg319VKBtMyCQhg8D/MDvd+9+tn2oNRmLHQUpPayp9bFlfWv7JHT
bAsL4ea9sQ957tf5CF0JaYd3gEUIrz2GiEbaKPpkXdBpA5IRVujEhpTkJG+VOWUU7byvll4zkzz/
fyhzXxv3vuww///2fvQIelJUnj6APZWyPKPS/GpON1BLbfVo7jZX/JjFAncz+R+EQMkI1LYM/NtZ
wCJ4jAm3foYPyIh+pgKWq3ZEU59EenoI7WNHi2aY400pPTFMGwD6LGChSO0DbaFcpS7JQMCMrnG0
QBSyejNjNH8gZZF8oKAL/+fuNjAfHOPh/bJhaMMuOY4T/EJYnJYf4HMgj3CtbaGSFQGiIgHWqoE2
Pd/E8uCENSsuAmHJVPrJN4DhdSVVdfUbvqFsjmmVdqJaufw2jPF7uQyEbOxqbUdOiXgZ2aDkdwY4
w6hHQzUoNXnSULbisEiloJlcz8cXthchSFHaiFmg5LPGYbZU7muOTEUbV7jYyG4g4+t8KKgDE3Vp
bNupiGe2h7lJo/GRyI99XYCR0vK2c3gcnDSdXyM5GKSLz8zRyjNyfFHkRdITXhzh3vNnp5ynnzx8
wlD1zo58WVb9MhQZm7alVa1a91vY74/J+o6VrqDaaWWS1E3xa9t5crz1ZNY5hO8d/gVEgAcX34x0
kuXRMPeIo2Cq1ALF1D8mVRKbuinINRqxVC7fwrF02cgHTK2xvIRlVaYolRwOx/WTiFIrjsxwVrJL
Wi27918FKZ4kadeLjiReq5ZT3Z9SHQUT8KkfoX6eCs7fGuqvXJ0nNRCzlr3nlaPATkpCSObYJ3C0
4oJbIwOvV9ed/EHVySeGQL4d7wMOIbBpSfP8r2ZSorzVnVZB9E92PtLE+ujggz469eP8i+NVZfnh
obFp9axMsAHhL5+V1G1rXsp+4lFcpUGx9mWwQ7FMfk5c20Pq8ZdVdDBOhYl644+KTwkKZ95SU8av
EKQLirlkLqdLwqrQpyKsTk1RKuYVEznYvUbWcftB68XvyDkqnp3pzoZ0tM2xiTXW2G//ArSJZex3
DLIS8TTgFvwgG3i2jjm4KxmLF2U+FLIZfMAjLDYUmJxxbn29mVbYwrilI7JdEoY0vE3Emc+RLarF
raMljwJDB1gHybMuK4PXBSHOxhlvCTdZhNzGm2WBKUbbANXu6BN5WKeFSmNspnIj9roVvt1BAu65
3ECXSU+O/3HvUqUl5T1NzF1OFKMXgH+46vs8ilzdveN5UGGoZazbyskNwtoUsOiXi8wKnsanP/7E
K/J3cwql6WVxVhHd9gvT+w9iWclmmQsddfahrvfE28FVTm8QBAsP0bZK8Sui9xbtzg/q6Y40Cr0D
c2ShsCqHIk0hU7M+njDMT9ufQsh7/EbZHZjNqIb/nzNduzkHwkxgUiV+hohLZtVClB0swtleh4ex
qLMN4YYH47c3g0YkavaAHtLHpECpfmD/3s7rhcX3KIyBAScrjU7sANf2LxPDcOEyIv+VRwdcApYF
sZypeRWjkcIzc6B6NlEsPDcw9dW8CiXt1dOIcuZ95ETuCeGiO/qkmuphrCkgX1kOQGz93HLJ/j7e
PjmRx2tGyggqRQWSRkgbYaAGkai3khLuPGGk1/t0P+0zGjwu6VSty7E1SMuqvpwJahRvENh32v90
m5qp7ioVap8iHW79Hnt3Qphv/sBBon4+7ZfKAjlm5Ij1LZc0fkVYLwnFHz8KhyUVCcQR+/UM3z+S
pkAyImTY2MFfDSkYMUAbJWHU7vjLNTch+ejg8cZzceDqeT/8q93pbyL+gQLIrOiLRr5gzjnMR/6L
6bGvPPZRVhRekdnlsFf8O1iQO2KymqoTUXIIVCEauS+mx3h66TUsWF1qukBHNxqu+Z8C37n4FQvR
onIFZVddJyspA1W49fq/gOan2wKeIRLQmjY6rO2Rm1ej3qmFX0f2kZ7H4H86pnF5ji2vrJXqkamL
f8tvBWfX4cTEOdvqT1PBccVfgfxUjOExZlVkch+Q6COrN6QGIQ9YFVlAzssDd1hGjke9FXNSP//W
QQgBt/Ankdbow7yePixaVZrj0dOuH8Kn+ipPDF7eCJzYKU++9b5Lmc6iaXVFwmgm0Nw6xtg8SK2U
Iz2kn9eJtb6v4nRMnzwE6k+I9KXyNr29++vQltImQw1kor1o/2Nn50vkQG0ar7EoXE/y7m89hELJ
Uhb/jAXO7DJPVLn2tmHyFm4pPFLq/IREk1ri5KwsO5kUaCbWMYOW5i8NqB27osnXK7E1y0hotepB
9pSjL8+18w3rGrKVOswwpczRgnAaD92ef1lRslKcTcKFD5tQrmbpWEXP8kaBaCBw3x9o8GbcLOqR
rzIx4FYDz2eZgfxbBzg9I8T764JxIY48VnJgCxGWrPlGha7R+Ktc/C62f7UyuBWcIoQ74vwzGCRz
wBrAziaYI1WzNXW3Qe+mBOoXH0OotW2ftYKRczwtfGgDxa0XrjDmb05Uk4yzGECI24wHXACjcEs2
i/Kr5QcpOUYNlcl7kaYw1Fak5M84x9OrL+GkASoxudYBoBJNJzGCzJxPTxBFxB3kM+L1mK6A/oIW
EAJx0Ahu8ofzlU65u3ev039rXGEm20VobHQShyuZ+VRJKhJIcysy46p8ezT3b4Xgju+u1B2RzfJj
bKphjMq1663uhLXjzqlGMc5LYgdSBjQLeMxh9hUHx/MKFOH/M6Zkz8wNULrxpcD497U6lpXU9oxm
bWQKANpw/CxXQs8+ssRFCy73qJdvlyjC67xaJaULb2nFVPPm5vFurE+Y/Q6hg3NSrkFDumPWP49c
Iz46HhCnGsBQ79aW9Qqh6cnaF41LJal7s1NqFFW2srAM++2jb8v8DTZNa7d26yj3pkF91NB7UL35
Cnm0p0QFemxROgxIOtVT93Jg2CO2Sn5Fa5Xvtk0wZRkTj99AI6lXtxl4qGU7tki9vaMn0pw6ROW6
5FUF3LJo5l+xnEhwC2AQC0NB6Bf4a5YauC9ki4rBoP9wyntf2n3NvPuOfRXvXR/BLPm8toB6UEQ4
03cFuoyGH5akqfMQB+tU+asn9W1BoHvoXzW7RAT+h3MAERC7Qi/V7Pv4iLJC7IMzuYN3VhFV5x+d
vobvCGjezbMXq2MYEBqy27vcVzeV2fUeQqW7gtcSu684yowbeqkE6hK8/KTmD9MLiM95jRBa1sqC
b9ozH97M4M06ER20AgeBYoRchyur6Koh9P84ccfJcDJIDAgmfZNZmkiX1c8KUG7fSZR5BdHacIht
kfRCBlLvArdtkF1VCWNFFfL5Gvu1HV66kf1zJtRGKNYdUV3ugRyXO1H3ubYN3LPs34P6COTmYoBa
0jp17dxszvavF0IbUrzBVRE6FP7Wt7S9Ef3ZNTTk1Rx+udy/hFSIpecQML226fSGUGoRzkAJS4+S
bqBCYJ9P0fEs04lTSzZkAfiiC7iHSgc/cObgigiLkrX7O8NlroCMNDmnz/s+5jniROSXvoBFdGfI
auoZMpUT4gCnu2kjSruDXRtaeHbwqaNMATugl0SxD/UoI1g5HbufbO7QbSOu/kdSRlzfBoNF1jYJ
2UUr5RYCf1P/N61/0ZlmN41sTW3j8H8JSm4/qhYwDPsXs1084s/BWjuM7dIs4oPlnETiAsqZ5+VB
nsbB8xPNA2QCn4e3ViXtwXyjwm1TfE9rmuIg3FXqNK6VHhgp42VvmhpNKpS1zUshyGfqVi5TFMwG
q3oUD3vyURBEexzRo0wm5V5RA+2eL3k+AMSKefk1LckUI9qvKGNCMnONoi1434oPP/QKJIlpoo3o
zEsdKYIR0AHRWWvideGZW7+tP4XSbaNfUn7BN86QHk6NKIgLljrj3S79AuYtqVMgY0tjK20lSUKF
4ZU7mf3tKOns/cJtiLIUAg2O275ziCYkAmNm3Om/2uu2wRJAd8+sonS9GjmjsXWzjkOVbtJpexZr
8RJrngPOYq2/oOzLraKY+9xhR9Nj6HySN6gLm+rl7sDW4rim6ocGhXOjjhoc0bLO+iEJP+GL+sEO
ejtC/pNN1iPjzxav5u2o3GamXLLfLNtaRTTDHAMsv7HCPpK1ryJneWHE91ufB9seYIC8MWkTz6Og
pN0rAUJoEIJYGsbz2j6e0JcKmN2iMp9AGbefHNS4A/KYnqOdwOzyrWoe32ln5zVLc6Eu6nsixUWc
nhF6afMKoiqGaXLQfRwEln6ve2zJBsBiAdSRiRHOrmNozzX8XEszdMa308f+tmVCytMWBR0bOXCh
32z+KjTPmIxfCvksPUBArgATYoXZU30oEVY4im265rfwFgG8sHG40iShXUN3CVoqaZLXcxNTe+p6
PjTUuAj9JORAkGiZb01FObosCeICR9qs1a16wWTmjiKtL8aHyLWkEaO8zdu2E51i+lGvQWYR1MUZ
P1rsURA8T7AUsPfjha68q7yrpO04BYqcpen6v7nImNEf972hmrKTW7VREZLWeD50398Idhsk/TGu
1xVxdeK0O+S7L4Rj7QNnVuq3XC5YIRyfqdYYQcOS1izbhbN2dT55M+Bozr+vk/rPk8lO/5TnyXoQ
O/f2gbYXoq+1mEIhU6WkINF4azTRgn8jVQFVklwdo8MxbllQXW3/MiSO8OD6UUOS1+uWCTweF/5P
ZNqwhGs43MlEzZtoCPxwQPItk8y/nxk86N0ggNpWEeGeC44t/zUB1ChApTXpo5udToVpE+odYU69
vIo6yPCndRSo9wMtrNQGywv1k3XZkQaG574yd4YhN2GmcoDDcap4FIUSREFo2GQNasaBfDdBSiGL
KCNj8ig+hxnEeNeJeinNGJghnpQG8q1PHmWbe0dQka65JGChN3a2liyoqCr8Nbd2toqcHSDJqjVd
FHrjV47Ud+ua3sxURd86hGj6GFge1laiqZl/vg9WE207eDWnMlXkxMLgdn/m6oei+f5lgB3D+qj0
xqT/XTuM7SQ6LrZD5cQbTHi4ssJsS8ZafxOkIDVfZdwhm1vI9g6ewAThlVXqVZOYlD5Ab+A6MuNK
ZyAHIJUKodvdajoKUj01Ile3t11qFID3jez2l2s2TOmI+Q91wnYwGKRlKAotyC0kresotQZJN8Nv
hQBUlhgbCRC6ULvAUhMs/tvmETVNhvm13gXI9lZLlurrRld/ERi3aogbMc2jTMP96a9+/c/PjQ9s
6eTNX4Gnlqj14O7RJSdWOC7RREBCUXs2zLP7M8IMG9kfwuMSzsiThvaKgUe3FsWpv2GZnf8LAAEb
NoxSVKGMqQg90Kf6hUZko7XXyZ0nS+bLoiFQmou64C9fwgN7u9GOuuZ3SA5KSNwzYWHcCPR75nhz
9Ti1zJkGBe0m+sMGxH7/nrz1bx0SbJnagClQ2lgJVagwrln5124BADjcQ9r2NeYKzT+EbgJK75Ej
rOVgzhBXNrmPFjiEAxiRKEG8mNu/dgYO3QeXPv9xAjYZEBaznWEQJa/2ZajL9ZaP04ZubFeGiGhk
r34PvHPZPUfQJBcvKkt+fA0VOZ2zn9xaPd6yMSSzCs8raMGncwM2ztOQK1HwYinSWwCuPelwyY2b
SqecOVHC6g6psImnxFRaqc8yG9priQCqfDSa9LsNZTfNBacOdMyM4BFZ2lvUsFj4wNZn3Qo0gZ7X
6f8U99T5ILzMHzT5spzLoCJH8h0HMiJXlkWwtzz1rn4UM/NJFyt0Ol4H20MGuKwRQp1BtmheVwic
CG7MavJjBMQmI3sSgGFr/1j4aD6yw3twirFl8P2vPBg3Q1ULeWT6XjQdrDhWx5xI5sEFoBw5Hd7Q
yH5cCPjn8zdX9/JlFElj7JW340JABejpyr5fhz31/PTM2gXPu3cvV6VwjDkXk8s6I9gLG5pTv+P+
t39zI9ut4gHdcgVuVnI5iOvfazQp0i2rUM3ctscPmisiCnNR+CJELsyYPK/sJRLpEcdbAAiQUiRJ
vOlb08rnQJkL2I5ku+HPtTi3vvZDMOFNqDC/udo4POODWKoldbsNfinuh4FB8px2aZ7i5rSD6R5B
9h7CxY0WLqyDgTFGSje/kMKRrqsEmEK36WxpFFVAXCTJPLthFZqLXkF3DE8n7xt7oQWdsTEDSdwY
xcu1zc9qcOZspskWeA0pK14Eu4WpR2n76jFbhO4NdQpIdJYpPnmYilAKXNkrE6jAAMntGYkSJsmc
H5Q7wAbxiSqfL4+aXLY9bPcB2Py7p0QCfcF/mU0Y2LGlZBriWpHr14aknrqm6b/f1E+LUhryKWQT
G9k/i3oBfjMKfnrhIRzq3M2rJ4WieGpBx0AbwVJE36Vdl5G6eVYZ117gcCUfve5cl+unlmWHz31X
L1DiN3UtycRvNGrV1gdJOD/ty/mUceOc7IJWy0+DijNu7A+1uhDwBFRn+5gxvH+PkL2gTNEZYtwv
yf1c8tog+7AXJL8SC6nbbg5fbmRFsMgZe0qomUxRcYI/rqUtRHAaIW+ZKdsPDGYDI9R1kPyhs+k2
UcwxjI3IjdyG6TyxxSrm+Or2IT4qeEjpg9shUMCAH6Sy4/3DVwXZAZehhf5ItKZ0PjJrDdOU6eDA
gt7i8iFys83mxqtmJYUGI7hrsZLBm1uKVK39miFuJLAkcdEudqE5yuSfnOM03plvnK7jUx5SUPtc
5SDh/ziJfAc44/DugcN9yGcjYqdvbdXzLLXY2CwphMkPRzqNC34HT+qb/KAkuiw4Fk7w7dHyIO1C
IDxij2I03aNI8J6vx6ewqZbJQTcJ2/3vnvV3Ui496EddBihHuJ+snpjuolepS78WKE47udjqZf3V
Cmni1CAd3TuxqzADzv+8jJhe1QT36XDDK5H1etWd7b9yq8ZHPJT+3Zwdb/hsRlQ73BlEt2NsohCl
SpZ+RHpW0CT3ka8fDooEAhU6Qv4LWJrRUoWlb2/2/ntd8V/i0k4rDoPhjdOaSQKUcy17D430F1yC
6M8RGyW/LMR9g33vBG08ZaPKEQLICK7rbgzxGakU9CoodWRONwBFEz0jXaeQAoHGvrL9e5N8iwKG
Fvtncv4/awldrsy1NIF5pXoXudOkXFAO5IClPlISys47CWbZdnam2kgSmkiZOCAjEvOnk9qwD8Ct
Lx3MHlxVHti83zJSiMoMVKId+O6FmYSjTzxxt6Acr8p7WTF/DiRrG1NfLAEtP/CAUE8TVEKc45IR
iOKpzKQHnK7LbxcvZpkili5oQnBkKSb6XcOXY4pNy2b3kHsVyHV1uRcfhGHyvGSHLx6CVDJX3Xzq
BG7AaVyzshrZTXCL7Rd5yg5xiEUvhJJcCk6l+pnY9BB9nn+cOQmdQ4cdoDSA9qcO/zBq3KHaPaoO
EAgfuH/+TgsLP8FRPJDBthSC/+VKW3TC8Yr+H2x46MxY55K8/dNRRFf+yCiRky9fePy461CjMziR
WG9HmIMP1Ufwm/0UrXrgg1bnfhtCfEXepOYCTS99RDHo/HRkMyQGvSdAzE6CaPQpLuqC2iYogtYT
MhwdZb+pfhvix+rycn/WU4TX5qB3nIAEZC/ra5Y9Mo9D3n8XE9cNkKKs9o89D2UuhS8y9Xt4Y6XK
uZlBSAAlAHpjFP2WBPmaFBgk9r1Um0jCbHCifU9rTUKDbrl8yE5IA2vgZSPMrX6VxwnnxYsK6pFs
Ei+fZdEGMMjntH0gI/XBGPWoA2c4Eve6Px1xm/zrys5iH27t8jDW9zXQvtGBdQeB9Ht1N/qSp/r4
a1jJ8IO5PJuXpTRyhuiyMFRAFohgZfbjbEeNIfnVX1viVDOL3LszpZ508cSvMUYNPU4E7ZrEd6iq
hlKntWm2SSSD34bYt3GtyqAo3Q7AR6E4Ib/OctwNOO/ISujLXIBHVSj/KEghymivhDZQPXfzKDXv
1WDrAw8L4X5B2T+zVpH+c0bI46AhwOGOI/mMLQHbcG37cdeC68H7SZVDnHmKBhKirAKgDnL16fVO
nsGxZ1tXTFp2VnKrpLZ+JMi+Qdf9gwBSyHE7X3RZu+N1eBPbt6W+T1jI8lQKChaYs3AB2TymANsv
1UY0TuKDi8kGMIkrcKRhnWyGrK8PTmbWSKxagKwm2h5jVxeZvNN19Ql5MMa7jp+lwV1yIgsRgIWd
rbhzBwb/IBb7MiTRbbsW0FehQlaLCBVYZDjjPLnFAbxE4WR9Ffalh5yUrCOWP0Hem7l3bRiP8yBk
lB+cFkCKwpA7JtkN2odlcEczhRE/NtN01xfJ4Ie8eDClYWngYywrvCe6z8xMCchMoIg4IaMuIZqU
atQHXHXnMmNUrQ0amtPw0/ZHxPox7sSwLMGd/CljxeaCipRMhoE9R//QZS6f9PyxpBejcUo58DdT
s424QU/8gZLWhZvnFPlvdQPp31jnEJRmWFCZGgieMy7tYa8TCf7JkkyYsf1d0F+Nxiu0QiH/Ym0Q
4Qor+kIpust6Cu4Q4qTXY8BkKFLKsEjtC/tBDVJBoEYa7D1ln4hZPemmqDvbQYKkdffcgJ5QbIst
mvnsdHK3CaJLWwaaSbznU4s8xmYODsYSD9y+umgGmRW6kLQYiOuJc5cPGGA5rYWMuj5O8cFGRBgG
tY03ZAUrYLoINlf6J6WUEvb3UbIJp//5kSCS28Kn1DbOFe3S4Lg3xlMCNMpZBRe/raMr93UuRFtQ
CGy783+NKCXPWNxgb4+/62mo6EeEWliZ4z3Dke1A+QlzmWVHjmaRA+1FHV8mC18ZrxiPPi2Ez+Dd
2eBOUqG+LmjRJ2uWZWs7QNWnK2fIvahOT3rihqEgQCndqXY60se2NM2Eu3IaxFy7rZV0j+y0pdbk
iurcyvhV3Ha52VnC4jXIKZwwKgeRb9KKpOX9l/sPImMDNt0oeZ5yOs/y2LPAIB8wfkSs0oIJayAy
RwRCH9ZfuQrGa0Ts4Voy/wXx1YhE6TeHThZoF9pPw3Z3+XVJQVlcup4d/vArvRmj1UcoUb10KQkE
iaw/V59Wh41oOq1Jv7+D/w7DagRYOgwePAajVEAiekXnVypB47r6TdUsPHVg7JaH53JrPKDqPXwo
a8po7mn00/KJNtoNmfR7pOLZFFBgSNy55urHRuqwYcaXp32XcmBbEK28ObvZ4SGzY5UxFtyJ9Ye7
xtNGRQS4cBfgZt8K1LxnTS08xjWcK1RzPYZo8Fc/Kcx1ryLSlqFN1RrMJYIBSbLLxqgutI330k02
1SiOKmkf6SfDbVJATGvqZHWJefNJ2u/2JjTZ3BJdayDJBJliQJT3s1SdQ/ypCF+exW6yRsZ8OI/e
nsrxKgWFAZZYjFMFT8ZpkYGgmjJsExeCWpVrsI5ISYwrwc8+bjgW2Mx7APv8bp+KYgivc1tiUkwp
zfviQuzO8eQO6usERGSxW8ThQS72G9ad0vlx1QpK+HcZ4rgToccSfS+0d0UrbKFePJPCTyeWn/sL
N+Y7fP6deX+YF4VIIbl4Edj1eBtXdqARvmCFrRUpNJ2kPb24uGZDAnmmhNbkm6pQeBj64Ofdmuin
+D855B8fBr0aMU7T7xE4TIdbNULqlKqOj3bEJjCcsKuFusj1xZJ+k9iE52GT9tGb+AJ9mjDXAqSX
jCRq3w9dIeqicTEviCCqwnHjR2Yeok7vnEy4YaZgTyN0Nc+OB3a7w2JG8wyUIKNMu1bbjf1zINSN
Rzfkxmg7Np9DAIz/9LrVuKW2qxkaksIhxTyIkOeHJ9PP0nfq0LyfYxT96ALQ8MkFgvhp2P/O8kr5
Y55AYmqTjNMS5CGPHW/Z4laZBjgFp8iKh1PpOpovirkddbyjd4EsxfEm18n/3/yPUIsk5G1g+2cf
tuJLI4k/weNsxiZXuRICV3X86K6LnFSAJwCFNkqZqCJ93PhTyglWjZH8pixBLY9oWPmOrq6um2aW
I2neX0B/4iR6Ag7XFFelX61rm7xBVrDLB645ZYpcS/oEEExh31/3TXJdw1EfORyqVdWl2rukkAXf
XLvEUHV7/fCCiX+CD538MkKNo/IQAozFpFCt1dNjWw0ahIXutk3t3+/BOvzPS+9EF/6Ha5xQMBkg
TrvQ+2+Gt9tkrRZvg8Ozwvi9mcJpHzA3Xp/rGzU4yxCedGey+l2OJuTgsPAE6EA030V3g4/c2U/f
hFsX9n3j4e9OD4tlI/qLWZJPVHJCmt74EuKFCJ10vjoeuMNpoB0zZbmhenGiaSBjJdi6/MdP8q1r
CM8973V6tHmLR9SlpBjLgdX8tdkxEs0EnDmMD1iqXN7YwnHjIQW3AOMCKxYJ0Gex7SENJ6wI4Obm
wrrjOnRPTAHn3nPDVRVDUviHPzJp96M3jiBzMLFdkWqkbWV92U7dYvSrxWak2smgzr+tEW5pleTp
D99B2SccXMBUaU92zdMUd2qyCE1m5UWZ2In1lt2SEH8XoFIuvxW3HJs7SIv8M4Jft0BNp2BmhRVH
jLrUWdPHWFW0LHhWuufASltKwBFXh6pFWej2GjmkxMsCTTaqNSi6oXpRDhj654m/wbNGwPJRGViS
d4+kSj4aCQe7yI0F7hmmxQy/7bwr5jqo25xrAYukMWWkPpkG/9vw3E7wE7XvPVwh+rw/eXtqTFAv
xXvMwn1escB0Kcskepfoq5Uo+azw09o1qB42IuSjvXJOFjha2cvMlWSXnDG9W8BJAvZCG6Khi5Xg
eJz+HPP7AUNXY6BGXNjfMwxRk16XR8uV6ErAmGF6WGrSVTtPZpDWejOccxpLlF02eLP53E1vCtB2
dVWmshoR11TFzsFRBPMJc4PyUrCeag5PFaW3++vv+9oD8OAVJiacZBm7GM4B/CgevNc8tlSgHkwj
xQlvDuZrnyUMiW2ulDilO0zbHnV3781to8VPzooqRcrBUCIz8Hh7QaQvnOyb5LewqvUY9RU9JS3S
PBEwAfNbDqF9gwZYcgXSN8PevjYJl9/vGjqmjnam3pn1NgLImMm9P+rk7aktUeovEgmWSr5++0ZW
cQTRMt2u40BxcwWaIUzEhtRsBfK0k28MzMiLAayiE+HI5iybRPUjhCV2ddTSA2KxhIr9BsviGGQJ
8DoJ3y3Wy8Ts/rq+4+EzcMW7FUUbvKFLUhxkSLwhgPHXMBoVVIg3F6k/7I4eW04EGpNH/FF+NCHR
/IO4+rkwgfZUHLc2M9J1vP27qo5CAf+1Jvo94Gz7yHj2VKvVHs+nIN4uUAyj9vp+tYkvGp5Asd7D
P06RM6HI8ZQu+H+0zNBBVTnr+Y6IXp+L6KXsljGaCOVmlA5rQkslPLvcAQJs/tX+D0YOwEX8mY7i
9XGXh/GV9wsg9ODZMJU6zztWKO2Y2WHgUe6B6hdwpSfPM+VDLUjKKbpwik/3mYMqM9Fx3yqq1iCV
s4ih48J0CH4vB3rKAojFlzxx8w2RlufHJhZr0bCBgHx658nLQ+7r/MJzgIiOXfg1V7IufJN5tmh2
5SuTcvvEPuortuRrs9C7Rx4AAXN8aKYd8u/fR49BHUDPTCXboO6lHOUtLo3wJZxSHljNeQ6hTC+e
puW0HZJR8cUepikuBTxdKHSoyTN5nm9y0ks14872RLwiNrdkK+LWvsOd4VEeVYomBk0+zXzHr3HE
Iun7BH38BtfsuFOgtRL/pC0YvtjFE7q6CGsTwxyY385bEtkTdmgMbdbOeZmf26EuWwQ11yKlJslw
ZCrjGbDuHksbUV7tG6XpcAWYtUjq17MGzSEKerZieXeJPWuoxKu6rpB4UE95fD4juivBgQB7/PPP
kr1/SvNHk7D190M0G8CMiQ5bpJfnkYZJ6A+S9Q1/denOefptQeXVJNTZKo6NIPxKceLx2ewqv/Uq
YhR2bqgbbxfab9k3lMBYx7QuPS1UZmnw5nLBjn5nGeUe/3zvMIQqvacKUgIZBvl855AyrBQ/QPI3
OpKaaDesPBOF7scy5MZaYdJAVjhpvWk8QKZ+nyOW81C5KIt4r5gmsPDyZw2+hc1gePS6D55FJsVh
sUM8BWVF5QlxqG0nnvhb0qWZfcILnaW7C93dnAGo6bd4MkEeoHT95HJy52p5wW80EBftDlGZNDdK
WmWBK1O5xuRIg+sufepkSA9qP+QT7+C+KtguSVRq96OHVspSaz2zU+CPauHSnlAFsvamC1++X395
u/jMQlYVQnErWp74jkFIcL6HSum+0bRNS1d11YV3oxbAF2obflEhmGFwHcWS11oE3LCK+OMxq1pZ
UX70x/Pn813n3P5INzTvgXrubejS2WKIM9RsxkaVaISoAYRKmGd/sDfQ7Hc3ClVDOtAHZ7ov5Gah
2WXdCfo0Z+QL2kVXJ/Azo6wfvdFnryDma14mL9lNy6bsaaRSmCkD9aluc4oP9ZH1Rsig4M7KpHaT
PCGmcy9XBcG10uhxINvPmH7FDlCch6VCpdIR3XYkHEJHKPeCEvrBQSzoddBG9kE41v8ttMZbFv5Q
P6Tyxyp6K1RERNQoEu4bi847vEONjKwO/PIWWcuHlLfe+OWSEXfZM9bACHt5ZxiaBfls9p2qjOgU
6wzE7AosAAoj34WQb2WZXuC4HYJf4an6x/Z3b+hYgt+g99GcA3GdGjLQVS0eJk10uZDrTArqOr0r
cioXMX+8vKLrnhjlZ+XXvHFfLOL7QrwkmwSDTEKgjwMt3LaVRClTu6oDl2VJdwUfF3x86THm602m
sDnfoJY/+OVRi+bS5SHBoal0LnJmpdTUZY9X+RDlCqJf5nswKJumSobUdvRFFh4FWm3h6zpRCELZ
se+FfKajDL1PBvDGSTPoT1J7aH20Fzmo1NKf8G2pluhHJn1jZ1P521ENpxec00YoUmlmobajv47q
NMo1fYkN+VmeoXltd1Q5sQh8MWc0e/CzZJx/FX2fdyiO0J4KfFWPjakMCQynohJXTTcN3W3MDumQ
h26zXyjefdlUr7pdSs8vRV70C9eaLvQDxEqI5q+lISIOt9LXbhwtSs2TrxKrvjEXOrocl2R3XV1i
W/SdGEPQAqFaFlHoZ7TuTWjSQSsdfopnFcu92aSrTQ4eRR6JdcZwD6jKBvimJYiiekG4rFJyaDQg
n+x0zb607b7eqgDNtmpbTUUgbL6etT9yfb5g1LW4SWzYzUxydfGwHcC9IwlTGEIaV/Qu656pnCRH
MVIzkUewustHIRdKfuU56UMK0/X3OyL6uaNdYF44FNyhpfLR5eeAtkDKiRG5ojwO7dwC68z2d8co
yOBGCEz+Y0VlZM7498K5IsIR6TDJPGouVF/cdSAn0jGqgsh4KtKhS7HuCMYLSusabVtloB5t4qmO
vIcCzwy47flhM1UjT4waCvnqzMp/qr0YpQxdJWb5r0nZPvJ0NSiGguHydkoBKPwekuPk1Fp9LSEh
dJIYsU0gtHzEenJ6msKQtykWMeqe1mJeFdW0czFpjGyfjrK6QbDVkknq4O7RW5HctC1Rx0BfyWt3
j++Oqwf2VHvE6HGbhqbw9mzo/u9rMiMvtdVatYP+hl6tCliW6/S8sTv8yPtWaZj/9zo3u4cJDhMK
Yh2UGN2h9IhLJHYg+cTGfwLFPR2KFfSftJhYT/7RsUmmtd0kZBRxu4QZySX/5UL5lA4FXgz3IAOv
oAOQDiIrB2lXLspdhE/Yr/jPUH1myCMULHhqXXE1vkuP8mLgGMaci+KMNzOTP5ku3UQ/ehKfUZy+
F5X+p2vMhfnewfb5/PAOF3PM4EGH1oafsie/xTDDft7tP4QZXsTMaSXpteM5aurlawqszBEDFcIq
1Ck1V5oJ/O0pKUA6gX5HuZUkbjm0jY+kqUtO1zHTA3J0ewtxcA/aHvIrrjYyC7Xtb7oDo9YucuZ4
BdUZpvt/W2hPlSg2xJB5RHn07bmXznhfrqieM/ZpHqxLBoVbhUXvIgIno6Isr9ZItnAnYOPfQUBt
KLYknyvqKzoGqlWC+3CtTOPoHbc04tV3oW3R+cBweweXX9NxvMM9GpIZTJs9ap2u6+LPo7x0ovWk
6vtC7HnIU27eYnCzK+vJxcDSUQqo0kabTWy66D6NOnjeW31BQ/pXiOwPZPMO0RlvnTJml9ytxB+3
ZjQfBOw2zTk/f/zB6+g4BCrLUZqVgNoWA3AtcASWcAWOQ78FdkFk2JvmAe/5NKaNCzeKBVk07tL7
4rVxKBq3CBBbdU2Gd0Gt7sUFhyeRJE5A5kVOigPL3cJtmgmR4bx3mNhuejP1xLxUstep1XACbXOT
LS8zltsTWSj/apjun57A42z/8VbrOgAl5fOWmQmNd3ZurMJm2uiS/0Btt9Fdwto+MDYkDAN6Wzha
WHw89yUx8XliepTUOp7a5rxUEOsz62ZW5lOkCtNfv39uEL8Ig0C8/iqRcolKmW5at96hVXRQWmy8
iy2+TFTLO1CgB4p4sYwNQXb52SqQT/m1zWU5q+WnMap/KOBL2mQ1PBZLfs6CVnZtv7hkb5T7Hh/S
HURb2kX4IyehSwHUOm94IbS5VWnnWcx/MBK2DLzxb6ijntZVYfONs7QLEHgAy5D0HqjwseFzcqOQ
SA3yxZjBrfAWxyfYMP/sEkHWn4JLSQA/T5v3CTzhcH0w0ERcoHhBJgT5UaTa+V7uMPp3pgtnmNzX
cuovqcrVR8WE0zUs4U7uiGmJIbB3weZwQf5EqvfXsA1unpxRaOySp2/ImR3mijy6YJvwSWqmBUh7
CHJbRNUGZZ3B37Oi06pZ3daCXIcBwSKclJifQ4YDMT5VXVGsO5EeCE3Ey4dKRorguYp/vj+PlD+v
01i6lRwGLxCqolNYxLUkgSAHwqQgieT4Ae4hWLvcUAPZxUFQGrFMxNM9a0gU52H1C2f2wc8mHJJe
+E7CIuBBimq6OaJ054uph23kC9ZVT5GE8I9jasFaRIXDKXo5aPndUnHSnhxwWm4qS1B5nyBWFvP9
jP1W22ycyFU1JG1g2iwrFlC8eh00EbfYTsVBdifMECZZT7MWGkZ4IClVtEqjrGh62alZgTzOfWig
CL1gaw4VoHCJ+QbKe5R/Jl8bNVxUcHSNrGg1Y4zeH7mwSjYyDvft8fZt/ust+SR1SS3+x6iYuGrY
JwsJRlL+GhTOmPGsx24WzbF8UHAnbR/Ez+l2ooKXCvJ+iGMpMIfdtJoyK6tq1v1x2VvnzGGVkqLa
LH6DEcDK/jMisL9dq7ZCgBNTw0LjsX9MnXf9QeDCGEL/SKMJmBPuFfGgHVhcyq/ZiGa7iQYUI+Gq
/brHrU97VVupRMhAk6rkN4L6M2IenvoA0d6041d+0P0JYLB2Ke5I9G0AW1OJEPbisjaZE+yE2vYd
uVl3jiiwzIw4EdBUCfXCB3v+203cZKG0Rq7k0nRRD29ClWHvyIMzW49VC3apeOIRbNU/vLe5IGfk
l0yWMhN+X6jLzlE3NhraxO0D87Le7gW9uhKZWsx+7P+bUJ5Csf+35wkUfp2cyKzyZbpl6VpZWiVp
yUeetIhjktvuZpEHangkbzbDx5IyHjcnyIcXQPaBncI6ayoMVyVh/6uwqcG1U8g6Ho7yUAkq3WEO
yxhe7YU73IuLfpvsJDcOpntRs0bmAxgFedtWFtZId7Z0vxSDBohx4cKjHuPmdfZ+9IdpIy/YZNF+
4eWKuXBjQBPMaGKEVwPGC+lkYx8GC9xSdlfjR2qtg2Y/VFex7tGlrEjg2Vw3g2Jij1Rc0NjrVqpo
vPuwWz9P4R5m58E5EKouO3w4f8npxGNS8IsbuLWAKzWnq8JTN/dZ+Zb7Ir6pOap/Lbr+ZYDliZz0
uWzstjOHV6aXZgM4fy1RJ7b9X6cwOQX9nHOzEdk9YYYSrhWoWXY4Fo9kfhec5U+m5Qjv4RnX7L0z
cef78DH1F0VloViWLrHBr24vgEKakUk5v/MYNcxAylE2PWyWOHr5ZcFhm1Rmk46iA+F7JBeQmi/E
blDXJUtbZyq9llF38uULNalV7jmoJpeZx3ZTvkHBgRCRTzUB9DMeSZdZpGt0tEeFWMSg/O74cVEH
m1t8GnfLCCPt2a4fIs4tufhtfKWwn7bvo1eQQt0zq0g47nhv28lmOg+N1uMoiqEMwBgx1dWO8fuG
dCBx8a5yw7Gg5+y1uUoh5lk8PP2tV9BgPFEa0lV7N77CXnIwyuUWrciorh3dtbGtzDQNQrOIGW6R
iJJ4vKfwrW7Sm8tv+LCS8/BtxIKjSgqQexUypMFOQOHP/Pzr8ozwCqwnfrYD9YGiywVurm7mRopF
hMH27P/Z92RYDO94Ey4KvSaF6Sgrf3haZAWe/IQL58Djy9Gk2RjbjVKVA0FmJrumbQ+mbm+KU4y5
cG7LsUcrPzX/ylF2RrkPTpHYG/ataGgvUfExoInljjk7OyIKAS22O8F5DTmGMnzrqKgtOINLs/vW
PV+M5Z1BkYnOtLaJZb2vUVh8ZTBx29Ykn0np4RZ7/iCyxcew7OGkCc81ToXMg4M0puehxqaEXmuZ
CZh9hZ8/CfGqA3ZUEjzi4gSCPUwZWVDH+CZqItFQqIcupDAX3HfxqjjVhSuMMLG8CNHOmV/RXdRB
XO7mpQVhBSE+pxLVzDWTtDr0JXMQYBkz1IJ7UrefBz1FBrtlhT1fmj/VGEU/a19xfYge7AAQ4ZUM
W7Zgk/EsQXQvGFbx4oRLbjwG2rp1OTsQv64JFaVYfTw+hXjpqwOFkVkkVA2ydnjoMuChVgJ1GbnR
MXZasKz1dxLXKpewCMuahaZhrQXB8inDbCtjQYN1RTXnQQpMrebZqkQB4Oep/SUkEAe3DoMoAeX4
2J0uOOZI4De/7rZWUDYG6w+D/q9IWX97IaOYlipXSYDSEKJy55hihNE5cV3I11osoMfR924a8lX7
/00NuTa/fX+NcWZqRUdyOsMjZ2EjTiXeJ7SHADNxgMNdo4i/DtHBp4npaxT9KMXupoDSc9exC+WB
a88OT34Fg8tD9QdUa2jQObxWi+OFHXRBsmcjFM1YQeIpOMcNS93kIS7lVpkR2oZBk0/VBFFJ2EZW
+gqnINJ8bL/zQcuZ9u1BwoPL/YXRBwqQ/uoWX/MQzTGT2wdvPxvw5QTnuKcPAB2lAkSV/byGFjxW
RaN/h6eoRwMeBByOcdD5NHFPsdAqsZXzA5nstCC0kR8pXVFU360Z3SVfMihG70dObkFavPC2ZUuV
cTiwt50+XnOTwYoGnLHdxv5i/X7/6ue+leXfgc92IEIyGXEYkunDWIcB+xV9+2w9sG1H8FWgWAsU
9zkl3VZude+4q4IildzNFYMZ+Ifrn/5sy5zYmLbnYOf0aTPMcto4ZdO8iw2bkx/+x3kzE/QYpjDW
jE5ryy1M/Y/dYsqlcbgXhcEFxoF4aJbOstUKLitUZ4yqPdYCglTzzaX6dVjISTZjoJ2NXY4gLTP1
RfaKG97sAwpt/ShN9g7V7dOcSYCUyGjNbh0hMtGgd7v8xCGzjPReTtyDQDPOyk97CDuJxGYTEqFv
6SOloBG55W6zJNf+zMaEKvv+N1M7h0+8ToKCl/MuauqHGpACz/eSCFYTfwZPZ69BW/Syt3FQDfDz
H/wwK2VfjXM55KId3F3FD2i6q8Pb97J8dMMfj0mt4orVolfb1iBzxI1qk8XI01nIOGbp9ilrwft1
js6A7IJH1a6JhIaMI95gRgOBebXA42i7r/OSH1IQ786N+PKQ0m+JRIZdC79B301oFmaS964vWgeA
bPI4GT9DYl3aBXZkrYu4dKJllfNbufFuhXWKSjOVAwgEi/Q22TRrYHSXb2qI3BUk3Ths0WmVfsk1
aPjbCzs+5LxSj2dTNufDvYYvai2hHSbSNok9oRGp5y2+sYc5vH/dOI0Ce3nkQWqG3kOCuGJQG1RK
riFpPrKg+DWdhTNymgPF4pRBfP6OZ/zF5GJeUdeatM6p/Ct6/NBxGzKW4W/B8zuwDf0+1ugKkY/T
nujfezkQu2KaeH5JNRwZIigZ7lillon4wFQxLOW5964hmdceoIHjCV9PB3THoUclc1tXTNsxO4Z0
iaOP18Id0zlZDHa4T5LEUG0Hj1LE4BdX5P8kUYdK3E2+aeWYBc9T3O5agd0k4Qiw1GV3KKN8tRtW
fCmZ+WilWiOBT0LgN0IsWvAy3H8twQc6+AYVI9yRuyiIRtdrX1MJl4fe5Q5YT1iQgFMh3ynBKC3e
VCOjnEIoll7tzhHt+qShoHhsdw2OnifEYwExRRN5AAIc1cv/2sZNrs2wmmMB4kVsK2DW9sCZ8Xtv
bA912DfAG0GYrDpR+egffw/IxgTInkyncav5lv3oLMwzEZeLWSZD3TcrM/3EjzHZht+R8MJKN2Rj
sgJQLr7jmUXSKpruF70jxq3zUV6+hUw3jeUYNF2T12dcDKTpIfQlrd9At24XFT9naqw3H6m0mJkC
lUh+DYWLKMLdhHGf0brKTpiZI5DUDjRdYpCwdMxrs7V8JSnGfCbVwbQAj8zGFll69tSnAuz/WIYy
MPMZM/vCrGLdiVHDMhyA9kR0fmPjhqfeOUE93QLsOwH1VAPrGWeRMaNBvwISbNHFYBPInjmp+Wnp
YHwGPHVbHbGjKwhucGR2QeiOXAU6XIqKGTCl1jm5Oz4KG3uiTQTfBVMJenjzQDkTptJPGM4P2r10
j/t+0eO0vEFEJG2HB6w5vLVim2d4N8Gza+WQZzpsLOa48MQk4KTBURJJZwf59fCe5VX113TwEFZj
X2K7AiqQL6bujbdz1SDrEzd49xJdzIkekh7opa0aMS+xZdkL6gLl7LtiE7orccWYupixn6QaIpdb
kZI32J47sNkVFyRBE29xdrt1foQH0lVP/TgWQ4xnwOXEXfQUJHkDPXWh/YFwVh0CMWG/6t7xM4RV
W/cfvUTNHdgiuFKX3RtXciwQxRuAunvwyFlT7LGulwZGha5T70vcIg+SIUke0V9rD3LJwFfpvWcj
PrpkoEBlap3pteK6oi5mkyaWyx6ijuji9YbKLs/lZUEJcF1e162PSWIRIsqgybwuC8zX8kQMot4A
WOm42wur6YqfRjTlwqOF3aJk6JMlC585B80EdZuokP4a/IOYLy0h9vilnAB452yVlgN26BGbjYrT
uHh5Fj94wnLIOdbq4H4opfA80Ewz+1W3qJytewkyEHC8lXyDH1Hqw1Usc/ovtO9Y21bbatrfW56B
OBCsQlYDNo++hsAfjHs5RPMnTaSXBAuqDkzyHn5fsOyHD2t0KPsp9omP7Dz30jsKFcczYcBvRjz6
4IlPZWc6Ev6ubm9goEuxBqMHLe5mmVs7H86UeQ4GkvkY23wL26y9dYK6RnQCMLPYjdSsOm/pIobZ
A3NpYqQFn6yHMqs3ifb5Jcw6OjfuPuxhaLVlko4IpQHshjH+7K0vmvmsxjgnST3SMdNfE0Dmj4F7
taousg5J0nMR6NcNt2KkwwH8wi1JaZaKkueOWtwCLMXYpM1I492ZI5H8qLT3S1bj7X0xOkQ6QSLV
iCQDtuZcL0IkLmHczHbYW2cBdzn8k8meGdzW3wgQEz/PdZGfaPV8NA9Mw/F3HNf2nKTaktSa60Ii
qTK7XmQWnIChnyTPGEhWPw42qRZNThwfPCDpqPi5Zr5E8b6x9bIH87wHK/nufUSUnTll9grgoo2L
zMAGyJ+Ib39CY+xj0HowF8Ss2aw8bGI8HzrH4k7Em4DDutbb0A0ZDfIsi99ZjVcUDcbG4+h6wjca
Kg26kF6LGkS85961JiWV/227yFFoHSkgAmVMm8S9+8FWeRwRj3l8VSkEmAsB+cj9szOm7M6oe9CO
LsIIKKt1xAapP60uoaqy0fKJkNDCaem300aCqJif7/9XU7i2VmIKdIK3uU0+GFu4nJYodFpnz2uN
KCa1VwA9pFbXFReVUOFKVSsj696n5MhNIEIH2vQ0vF+3CgqslZV8DixZHNwx2eWP/7MMmMJw0Md+
bGhqk6W0YGDx3HFXhIbkCGPfmaRh+iGOxbqaF7O8qIOswltkTUCFpBUqGpdpFcyx9uQ594uCqIX1
S/c+dEh9MDIksAofmI2B2GNv3o8TerqaCSgDyQVXhmtDY/u4s0Peia6Xy0FkyitbpoNYKSqPUqXK
3CZjKX6elPCqO5LSkVVnG2tjPVVqpAcvO6nA6gjLEq8GdwSTjUXvDgg4mE6EvJF3GFF1qRZqsWoc
IzzhjkqyoveqQ9OOr3ggpjTQKnEeQrP2JAvmwyihRk62sR+BeFZidGdIMlO5zTeqOtcPzgjjnNg6
UzF0JwdMdgsH9PKLGG7kvtGSG3cwB8jiSClUQZOSMcAfPBgPdQPat6LKGcXAq4hllAp7hIRBen0J
Hxj13Ehyyvoy+WWrKI0i2dn9zh7VxIx2eFMll6A2jyi7jjOl+viHr6syyHFCpgV88bSe3gjnlvOq
Mcf9KHGQMb0JzFI/CJPUYW2FGZXGmoTtgWnrW5mZGK5nGncLZtQ7jXs58L96J02/scUZovCpP4PP
/ZnS1sSBxHCKs5hmPRtxGn6i54R9ET5f5XO8HY5Hyuj+smDRDJCDzVJqbdP8l6AAkJrj4PPOzNM/
FSDR7kRtbIxDs6kBOmzCL1syLiCivrO8wKdJ6aDduIEGUuJ7OuajbCkTM1yO8KBzqWwTN/Nt2CGH
+qhrZAR9ZcFOp6o7uTKD3ocw9GfRtCNvf3W/eiV3QLSWPfYwkrIKLmc4ugJpCPsJmo0A53BiZQWo
we7BEX1XTBNyDw793infIz7w6Tot4DGBIahyAn3XCnOmONz41xSh/hFFjq/In0dRGiOCOn6zPJjo
lrZHMcSxmhoxZzMUIrXmt4GKi0eyqY770pXQmEyV4p2t5ul5/aJSkmmQ2CWE+waGlv/Ae9RGkbUW
mvYjDGuIlwpcpHPzDslsqUJ06Iw32Lh/mxo4H2Jr7HXIA3yMVTKgw37eJcBDjXjU7MJPijYpvGCw
ijoVjQH3b/iH/Qv6/8XKx70AsTe45jDIEBnkPoydGeFywzWG/shz7PpgAUabgfWtXsVfwtbKYn7A
ufYRRfvkm8EwD4G8aTvYnqE/Qo72lOWyz/1yDMOE9jvqS2WwStBKz30jJHtOvY7U28PaDikSzOmm
b3D0F80xbxakg5n5j3qZo47vwq9DZSrFf89R21rlkNRvL+JJHdXJNiz4ZlkhphJvGOQkoBOTcKvD
QGFBRci4n/tamlzjst2TtyoHqihOeyGSs2zfRjFTo15KM0rtInaJAIfFUtQG7O3ijgvYe2xok4VR
NY1CFaaSOIJFyWTOvC96Yc2TcGVJipOZt5hNPkAU7kEDtSNSXcvDn9Jo3Av1a06635o0XzUGUpEL
ha//migmy/FHPRAmWQXSxs8R5nCytvQgagiqR3O2yVhmPPsMNrs7YZttPyqwWbvi1uUTTW4Eoq2N
e0gYbQdTr4QFX6X0u9cw+g928B/MvyBtkh36/1oJecmkwWZSSOF4ON0CAS8f1fAEDrxH8V69IyKt
9m1vAoahTMBsIiAbUXUQudsOswJD/Geq3Pwqs/U0ZQLerTzdvOuJ1hdhICDF0szMRrCD4RLVEgmE
Bo/kjNZ8YKA9Kii0av0rK8NgQAGeWicjrdiR7mTCTidinp2E+926SmeDeJYEm9kPX8n7LNulkRs3
kojaTuca8AtsfBCyz4d/I54OXU8Ecnp6Q9Ye9U67JYCkVkASxIH2oSyt71Zl9K/dmSjzMgkWbj33
oafKtrv6ogZ/OnksrkUXe7MdwCTdbneLJCvHz+lBNUR7Y9nFbocrppL42rSS+AMhzxrMUtrCpMnB
i9yMIBRRKj6Z0rZTmyU0MqGJDJ6rBAtJTXwGL9crP4SkBAN81zcG8TzkWazo9TjJSp6cgN1tc/oH
Hrg1TMfKsQWvt8Dh7VWEpcppPgqeNNHtQVm8+kMJ5Yunah7OWeyqJEQvf4n2opJLMP98pLQcrxrK
JT5QGyPQBbY6cRFxGr9WCo1+u0TrWJEvRB5jcDzojYXvSij1TtAiEQicUQvUW+mkvG4NNwWoXw/X
4gKX+yvpvpoJyTNkKRSDIBjIFmYuilFBo9ROL9jxNvSa4l1AURsrc5u79bjPsThDu2xOywEfYw/a
A1vKKk/3WZHwG3pGPN8mh/Av58GMKbfsTPyhrdr3BJ1RMTgVWSa12v58mc/8bqYJT0rHeihIvoXZ
GDSid38+zNsk+GrU0b5VUyKnUXkFdbCwEs1xHmZFpCNdNJL6KJAPcIx2uk6WMIAOFytvqClYT7NU
eLXSEMAMk8RkCGar6wrZFRxUHmBsWiFHNv8t+TIM2cHgT9wMh2tRT5FunUuqERvU1sJwdbEDF+SE
77EcOvr6IXitOeUQqteB0odhaaw9XMNbMbcJhpPCvzjFky9lkA5CQMVVp9SduRJYwnnp0ymJHCwW
S1x6Aa9lNvYqR9F8R9ExRroS1qiXlBMZQw5wTOk7BEc24UAbUVTcu34GdV7DZyZfZRA7V3YqgVwZ
+EklDlFZ+7ZtNX+csw6vBpVxqphgJR9JtrBvNWyfSzz9MbsQWIlHaihWKoCyCMDxcC1Xvst4wYMs
Wa+WdgqWDqxNQRRf2cKevHOOPSeUCzudXEvQpxtsaCCTTRLNy1QKvlGLdtJ+NT5tdDy7YFOuU0R4
9cBhR2/YRNYZqsHEirI6KcyFlkydMwk95bb1ewu08yDoSlaQJz/rq8Au9/8JozgLnXVlQo69+MOy
V9yY+zCSIuzLqluUYD1mnoyr2KBvPd8w7exsKFUEAF5fm1RseQKywA+Ap5zulAAP729ky8HBqHuk
KRSNIJYb6eKGiXNFsIvx13PwSpkUetNm5Br5ISv0zneVE/laW6ZD4GzNiImG87CeafNgASDyuJOi
mlDk7eWlw2EkavMCXo/YEvQEqjuCxyZPNkGMLP3RIBetnxlj7DnzC+rGfJqwMc3QjqnbJOHTg/BD
HDq4Hhh1vrIKVifv8/hpEvftQNsL/rJWUwgPOdpWech8McZBvBoXOjV8Qm3Xlk0qBbnb7RKMmibd
o0RvvXP2IukiCC7a9dZPTTViw2mj0GidrtuGb4YAdEk9j2Tr06Q6C2Wq9e4ZzmcOrsyOvKdpSNJ2
o/xvbZ3tnC8UnKLgrHcqwg9bshhrysoJHb2P/ImLZmUhK9FaJnn6TDRWApewUdEleoyBgLqy2WDG
pkXBQgrrj+LXvOnSylA/h6VJK9UWcgM+YCkyCYCoA27vwXxQ560xVAHfX/0Eb9jnf1HqyGZvxSdN
XzK9d6N27GQ/q35vBtKQzXCtEesjf5Zc3UNvFzv+MjnXNGhiAaRHDGbXadmUl/1L76oCKsECRkk1
ga7oJFg6ZflzjL/xyfu9vZY6mT1aWUgKYANYQIndBurTQqFJxN/yWuN++FZrlH6B7Cl3Dkgdzp8C
jOMDaEj2zQvXdFqcvX+ars6MKjDLyjCbapMEz518fW14oMDXqAhqn5bg0/AKiZLGmGL+jxRC6p/F
22tmrfbuLDIvI3r1nvmuY65muRDrxkcxP7idQt5yHRWLv2Zd4vj9I2KQldzorqU7jxc59M6cFC/C
oJ9ZTiq2/VqHL8kX0kcXzHsTRQJ0ko5/5Gze3MUiXtOR/dss5FvmuMxUloqKMhFTcXLUwjbmV5xg
bJXLhhE3a8GX3bIdxEuZLSIWKKHdgpjY9lzs6pB9PBrLNUWjNwF0ySnkbZQBE3rvhrdHud5ul9RR
JgkQXulC1yIOnWbyuZ4QeqbMv1afG12phtRfGTdcu2j5Ey15o/I1sjyxfGFlaQPDTO2snFasnXMh
RbUohgwHJfH3a0hwLbk8FzgtUnwyIP60WSAUtEB8ilC5rPz2t4u+j9wmvKAIqGC8M6zRmEICgJe4
OTTdfDmW4VE8/haFh++ektFfWXfqmcs0QBEv7q8eQ2xOjZXhJBDRsy+Iub1gprJiBxRj1un4lLC0
ZKKYZG2BfiNYLUyNwpziHKk2+OSnhQyADn/X9qDS4/msSUhIrxMVRkvJnVfHIZaTu+n0hdsUot7+
YTWQWgpJLbI+XIjpFaw3mtC+w5p9wT+ZLxEQz+vv6nDpPQ+K1rpKZ24JCNUtbcM65BpmHx2/EJnF
JOVKxYykqQnF5+H7trCF0xGKQRssFqkar4ORw+CgqegsOrjEAIYOoygpZpcXwVDiRDE7YoSN459W
XdcpJPcjSHn9oRpObf6l1G+yLuN7Hi1VYtNED/QyW+wvlAq671b1ZCDZzFx7FYl7fYrjINXPfDqj
vS5ybw6ciTRdyVrUjqWNkrsHLMxWO1rwl4yyE02fuca8w6QQlAlbvfRR0YdFvgOXs2mHFTGboaAA
NymblHgjZPpq1tl+1xxdGS0b7XdEu4K5wPBbAo5NJ0QxuVhbvanU+Bb4krB+IUqyjifPaDNDqS9U
Rbe7tpsE+mYbztNOSiJ77Wg1nphQAclfvK0vWxNcMOSFTXmPd7OuBH7KfvHciL27BhNfHCeSUDuf
Y/2XwfqytSevOIiRU40U2ts2F6LjJ62TsSaTpvrygIxFk0WXYQP0F5h1ZnQdpyoKo6ErRcPUstkd
0rANF8Gw2P99/tDIUrSIQNIy9z1SusLH0lT43OtglwaeUMr5IzFne9K7LZz22SiHncKcADMwIKTz
z5OPUKo57B7gGzb9DMxxgfbz4vL9Wt5reelFPwDx5Wht2T53uncBiPw9yQyci3JFvgL5z4542Fj6
yK1puh0RDc7h+Utnxzzr/cc2Ho7MF1tgqUFmjYKtRqDnAqZFN3gpZBVcuxwm8vx7/1cnkyD7EgwW
mwv/TQJQM36u0K5EwPOF74Dk4MZlKNCLQUgp2blNZycz2td4Y5jAnbMI4TY44IIjPOD/WGeJPRmy
JbjwPZTYmbYrp4p4AugywBtXXWv5RtgSSZJSdNCKHGN9cxEKFEGT7evlRZ86Q5tp10w5CJTS/KyB
BHiNL8df0/6UxN4J3FXDBUJgBR66Zfzb7irQNTLbeI9FEVpBTRa2UESE1yKvzawb32FUCCuuCl6w
G1e/qxcRkeVgrVlTXnyZZgfgVLny8LuqyMga6ZqWRhmhOHR5NsOeKB+vYIMS4lyvLza0k1ZJ/okk
qZyZkIFOG7dQaV/Fe65DOQ98t3pJvW2sYUx2VJ0yvxfH2TH0rYS481CcLtCQJ3LEqbMS75R/GBsE
KwPxnQzVbcG+/0IKPZtIJVaCJ7NH8QXE61ZmuJxc8oE6OTM0ycpvBMRpZ7EvQM5vt41nGpTHc0jP
T1PCBIGz/B4qrdA4Qp6ysuD9uTHAQoZ0jTtPwucRK+m3+qbfgpVJEGK6dt+hKWcKNBbkYlz3E+5i
/pHBRjPPhnnQTV8vkHV4HOMHfwsWnU/Tr7KlyxHG8ZqnBWxUeLKZw9cuoJWh1H8tgorvBc7kPYTh
l4vodKrVnorL0MIJcbiqB9C3Lp9/07mLuWfp5K/P7gVpQhhVcNU8bh5DRyN1fWS9ysRu0hDa5Ul/
/dhOXED/41b3cZPwp+5uHbOrMSsky8GWVIC/tHRtD3nFY4DwqRyvWevBX1u9Tvqhh4iHIYtUer1m
nav/uxnl6Dx3niYJQ5f3OThcJPRCYqryRe1TKhdhWk3rs1xoMmmpWjDokR3U6svNMYl2+GS4GAQu
EyQWm0tGxT0G8Y3BSJCTGTt2zzyStZnXQOQQ8iFOpic9Hm9muclRa6/q8Yyj+iGMAmN7FcJCQMWH
t9i80SBS/mtIJwLfV9rrgMOQfxsfUUc/xZkiQzqO1BZcCS5rd8TJ2HtRW3hnz1pE/s8Vk20XxzCu
GRSiwSMzG8qYxIAg+RpSX9h6Y6O3vm+SNKPyeXpFKjMrbdw+IHOznKzvnGj3dklfMr77mUzXqr5P
B32gOJt8LGo+m7xi7qSdbLSGWxAvlydijyOw2j/o8lVevaZhWt0+/x3/1IjusRbMgjhJUfqF76c7
LTUe+THhO8bhYP6gi/DlcsoYfMHMrjEOAsNgoOPg4M6dCd3JShu5eNCCjefpckAJf3iM3PNAFTQO
zlxW/Ecdu0xlOfBcaDHiY+xNKobWoCCdm7AEX/piTRVY3XGY8F3oJR8dDAE8HRm5HSMDa5l8pI8i
Pmk4xUeERUFtXPnHdqf5KBOtB8BjiaiyxqidY2pFOBNXI8g8REQdVgtLjaCQXUFmsrh5wVgD2ur0
uOOpqJV7+AX7HOzFjQnlpVlLvgTQaSeGjbDMVLIW5/kVo78YzinYQ8qpDYCf66OYpDofKAqBAosC
wd/eK42t8nAhBcMK9s/TValRiM+TdTnMFDz8GcsRP5Dir/aorRVbvly9Ny26A4pejInZTJV85dSP
0se+nWxHjLvUO2L3CAnot/hfVJXW+UF/z9pBDEMmrnOEfGYmMCBI03vwvUXwtgyWeIsHNonS2ZOx
/9xoIo8EQoSY+1erq/nyrA9CKDb7EFDcBNJ7iFWOQxGryxo3qHvsHzcnwmEdENif1u05LvzmmI5w
DcQDolmf9SeYl90cuZnUvXuGrgsgfQ9DG5VjrpXLAh3SjQl5+iAKmSwe+qpA2TrpsEJl1C6xN9R1
xwEQ7x36Ur5kLNQl5uV28pvTvK61a9wMVolNxPKNir+XWA5v3pLc3SVe/t6kljzwnmzqnRvIxzib
wdBo6bKZ/EljBAc0VBKmuQELTbHrDcKqf4UgaIhlZOvsx/h3vy4uvXHOaMsH5Ig2x9IsuiZ7sre6
2dMc0/EYsRDXuozWeVeziwAxYfkvnRMHMOZsrEN1ZTBqF/JDYzKNF63omPG0+I3XHWmhjzt3eAVC
vfrdJN1juWoJ4Y6a8VuuRQPEo+aGpiGM5z/C0l4Pz8yUpMaX1mU3rAVDJnH8DK54UwtvWPSX9u5j
awKoYnhY6Gpp0zLFAcXrH5W9wjVcW9C80YDDDNtYyh8DhmRto+Cv/XNIEIoASCZlpxZKb/qmyCgL
ighzhlqJM2A03py7Yd1PALj6tzkBZEsdgpLun2/e/7mJCa8h3H1FuXvBhPzlfvCimX10+85VVHug
kx+a5yfwvBYA6Drd9imPw8/tj+/cx/LQgHi8/gDXXLI/LtrieBQeWQbxzlKmo+ovud8uEziF0grU
gVUAc/W2yFtk4/R0Srxn2DrStf97JF4TFab8stvvWzOC0OaUunRaKl7hvRtYbuAyi1ct3Mcc/WO5
ySaRA/S6MXg0m+BwWqJwkTlpuUl6HbF+3F+i2QSSCzUn+v7V6QfOQQlVrEvvIfBwS0Aj+RWIOA1e
+WyaCXCMx1P0WrIqugiJoN2Z83ZqwsGJlpTH1VOlNkTsKClo9i1zWZtZKN2QmxFs77phFpO+nMPm
mDMHfYX8WhEjuJjtRHzznOrD/9tE/hcn5kpV0BN5tCGBxnVv7MpmUgXsNUxOwws8x8iHbvwg0J/i
564YgAJipeZuamA9MY9t75UjPjVY+uwymPxDYR5n8TS4dUoFmx4HG5tGb61g1JOAPcx0D0CUzwvC
sgRCJxvuqqlhKmCyr6vRmPUigBOksdq/SK3wmOZMM3ptnaJrIy7lxV+Rj8u5uBWRKrM1Hu008yBT
3vRafiKoXPW5mOssYfc9ii7UyKdjmzU3KSWkzFEMM2HUkuaXzE80R7kN+TDYZES09NPn6SrAh+7p
pL+4RS58ZwUpiRxWLM+zls0Ene9tclVBycKk5GWSR1h9zopFBrcnUJ6ZE9AUtpTARYZzxejoqqg9
3i0Ew3hIJSk4b7VZ5BNxfND3m1ys6RKbQqAocB2VunVEyOaAPDFE2aeXZhhngg4/ILWjgNvbjiWz
Xj2h3z6gS9xMAPdWNnpHBIj13o7MZhtH/3eZ1HvH/L3fgejV4kCDpWyZWDoiIMbEgBtQTSX1TMf6
Vj6o7TRC4Jse+/JeOGe+bJ9gXu+XDXVVjuMssz7rhOhQRIE6OboPLTvoIJNflCAqNv2rO7xWt3Fk
m3Et3Kj2fAdDWMEbE0+o/df0agM3FnmRy9oRaA3iHrlNoVr8dj9ZHba8C31kR8Y2ZyXDYz7wekuY
iN/SraKuaOgWt6d5kLk1ZllRahc+Lfn9wekiaKwJLxn81q4QlOaM90Dt9qpV0VVeIj7QQhhEYlT3
jdDvFoApMM7JkaBSsthxfufTD95/s4XUy/J1UkCnZJi3/APi2N6P65QbYqKR4nraDP3TjLHO+zxU
r6a32Rb8XzHwCccnNw3zcnFI8kO16ir5zz6qQvZ5tO4FspECjeVNoM/cX7ww1OMtjKnC47A3ncd4
bCSzmLDq6CdbKqzjEoQp6A17Z2fnulNxaucJpKk+erv8CZQUfXvDQ+Cdm5ugvIidPg3JR4Yqnx+4
Kkjk88rLgYMVZlnb+RpQOjqbJy0WhbwuQcd0WTlRoDmFfTBmzo8kWgG7vKzqJErQplvDL7rpyg2a
mwY89Y1fd5zmBP3hsKQaqS/4Xt88/hUD+xZd0ntZseroJx9/QWJuqY8GK6XZt6n9shZ/zKinB6xr
iNgai8uSIdwhdKt28CHmoEg3Ea5lIgrXR079YDqp1FC5Sh/CoOKeeo3E8QknUYFO7lPq4ukJxlbS
mCOFKluCFdmqfJzEsed541KoMidZ2U04cuAaV4NI/uhlqMsskBpjLACkQEJ/7f9zmKMdw/3w9RTv
eepia11ArkC/snvMRQvKfcJXBiqLYwEsS7XbBfQGWnqBDTJe3DQfwUT6oth+KNrFDUovyav3HA14
l0iQKYizz5QYbOJVNHW6JzGX9stTrpNJPJwK6LFvnAGKm4d4wLLs9Y2k0qaooyQfD978UZR8Ip4x
ShdEI3ZYl4qpNp6oOlMKLpFG2CDWD46yMjI7Cnj3M9edAkAFyubCgn+rgSqfVFqGMjZyhhTKYqfx
8bn3FuQddKz0dmy2/LbKGKMxPV6IG/dmu+mPXpEhs8os6C7z9IQ2X3w7uqAzmjvCxT1kFSKJOHND
N5ZyOqGToFUZTQ26XjgqLOVxP99vlOAmi17S/kDWfTktJoZnwPvcKLpFx4XYp/2spTRV229/J4ok
VMMvp6pMlwU4d1BjcTKYyiK604wzkLnU3lkCS4CQm4nugEN/8279lYBpR27Sm5Rd4hTzQvTEspgN
DWM+VPbuXoOBuqwVhdHq9xy5bUiGweJDM14IFsl/86spayLy3HB19w85RuG857l1NY//zluGDHKP
gDMxw72wiFNAYuk+jrfOQdAlsEYeE4YN1UXFia9iT5/xT/Tiy+csJR0Kv9sVyG3pO4sTKxFN2jBv
ksXMP9M6bAer3TZT2z4qlNYYQvDvDGipXE+FoPC4l3Uu5kat/VsCuX/kZYjHel35uPFVvTg/n2ai
m/F68esFi84XGH3qn6f8Ao3yohoI+z5G+tS+Q5wVen+cvgMkaAM7Op2MvJ0cj/3qzgQMeGs1Vi8L
NZMm9QAQX6vHaJEfCZGyF+fiy+payl0J0JawvdlASHFnVeb++V0vUKrF3YAeh65B7lxyvBztrHCY
CxKeZieMF28/toGAjnieywk4WqXkS3k29hIcwXqOBbHn6jldTfC3w3PixQ5NovlXPZItF8J7pItR
266SRY7lIDEf5vcGmKEb+PyZjfwpkUBZ95sqL0faVdzs20pZLMuGxIKuT0WGuGuk+5kkfuBt7LrS
W3qOf2pUzugOSE+OzuICjhqMynBPUxveygpoAa4MiRLbuPPngyCMZSXALD8Dia3TwP5T8/5b6Af4
0LHXgxqnyXYTwmtuIOvpK1h/aL1n//lfmQA/HD9f6tOm7VdTKKKlkA7tj4b1Kd110NfLBMAvTHxB
XsA8GyVcp3QNdSroz7RdFb3RBerCbZyyNs0EUz17V2NEgc5PmgmHN4V0kPLr0DO0DXDUHTlxXNgE
51sYgY5Q7tAmUaKWz0+Iov76aNlJsvX75uSoS0jQH7l4tVCLvX9AEscAiCA7ZTviR6RzdECK0wfd
d/2ZwgG2/TE6TV/LhFIimpoV5C4VwavNvppMwDkiBoIwhJVYIqTBb5oYVTrQnl2diMKkW6tcVjIp
ZRVQ/8Y+wze+eCyj0r0ZD1MDC9aQZn72OypuJpnDvxiIVz076ep5WRrvlxkqpXd1JVnHdml+Gelu
KxNzbP0hvMkMFU3bqIe1kU1l3cAGW3Tp725yIUFlYa9kei6gISbXwOVpWDlqfFdGKrAc1qA1v8jP
U5OW86Cs1jmAX+eeg1dRFX/GZ8BRn6gOKGH7J2PsK5fWtqOgUW+OP7/CUZmHNfytacE7t3U/lskM
7Yepr7p8ItI3uRzHqLryMF8RPXqXhDEta4NpCqOYnCmEtgdlMS+JqlqVrAoJ9urfzH8qX1cCF73t
7DYMXAgO6p8wyo1QehbdOuyV+yMzYoFfMn1iL1oFONMPs/z5z5yiTbkwuSioWM9lKlp0K1w9IzQT
q5vbN9HnMLSktSsQ61pgohFUR4J9RyVU6Pu/LxGu9dOWx5H+rEYd4k06M+0Xhle3cmEp9RkRybfX
s7WWzu49iDMx7r3aYYtuKLZlERL3Qt88uZKgvxEMFC51j/pKBvsBIL21KQw3RyMIGB6irOn24sPd
xmXnlNpc2F2FCnV5xUok5ms4x998SKoJ6Qy2/cb/AXAKyQ9+Rd4bDvTOx0tCYbHk7ohRdUv6hv6T
MySCw7sLF2fz/1FThcBytIj5lFaVQAUedkPKbT0Q7TOW7nyR9e6R45mBhtYyiq09tNIzXc0on38F
8rNAnWV2sRuQT9y3M2CbMVF86cKVWunQDRTUxfzfKos45UDI/CzujaqhXGGc9TxN2ZjcXegK+E0A
F5OyrBMf3CpJLd/ApX7wA6RpxstA829tmeoo6eq6pZXZlZqiVTBYV6s4lz1ZLQKDlfdT7LotMm7n
BgcGFmcnZPGWx1S25cFA8d8Cpx0lRDPQVdjjZdfNspjAGKwtezDdQNGRgETKXnoRl4ch1EtjF9h1
WQzaahcFKHiF319euBr96x3pWa9XEHxQ059gRCwCUv6zeMT/rzLxaIt7SWLE12XJorss09f+ZDZZ
1ujZoRAU302SDHdK185fVp+eGxpc+0cDHKBkD8JjKmMRCoNxbyDRqjeFHYrILIFis4Hm7UGIUzbL
Lj/CpfiBfnSNMbuL8w8HQZZn/9wtvMyhbzfARjrJeSRXqayHFXaFvWyf+pZ8DVZnkRaD9dkGp3ge
m/0dSX9mtQmqDiILeln9Y9TEq7GzwlIoaI4zJ3LKDycQxJGvoZG0SNTDOld+WZDm1hF1XzLtG+kA
dhjg6fKZov9BR9CKGP+RaO2bwV3mWMgy4AwyVxgofc/FI26ufa3KkXPb8Si8yOZuXk+xcXJuS9M1
3zAxcs1EPDvVIL01fQY08XD6WgCLHM9LGakZlhCpp5eN8DRs6X2PLuRmKq+CcEp2Ns8Xa8N74CFl
R2jN7ZGqvVOfhx0hPLLDr1qs5gJae/lmK6knTqc1ijLzAphFo2qtg72J7yNDHGZME1cxfHXvISat
qZ4hpasreJQgvH/XFXYbEyseu+vsGHI=
`protect end_protected
