-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
JnBBcKmCo5+q05YN9t8G0tNxe2max6SgHBeBRpUH4ezJLN2MH7nFLUas4iLS/lDeFWbQCLXzXtGp
zgVLfhaVBJ/z/iNeIA/yaVmVKzCsMMh1ehAtYPpVIqTyTTk5y6RgX2XQ8m2QbphGejzCDLNLh22U
zLBv7XyrJ3oyEcap7C1QxWjb78oJlX0KunhyNb0uutc2n8K3Mth4gLIimds5ctXH0QAyE80qVmLv
W/UmkIcNT8Zla/e2cMEqoHQAmArFuePFJJpkW4zgrLvIEaDnqLy7Ak/9yhMy5Nd3Vr22SO4s3efW
MROF3YZH4UXj3KaJq3+eKQuI9bNZaPpinXBHbw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4528)
`protect data_block
EcIP4T1D+cR7iBR1Hyjgb0/Ba9TKsydq9fUjx9yJI2CKic5L7gIBUXdxiYogxbqbbVIBXoEfEBKB
oAUrpoTS0Z5AYQxKRFS0pGZthN/MXT9iImpJIYkueO3FAGxZrZ16UfKHEf3gpgUMh76iQagQvZs3
VsxVFH+aD3FXIyJdNfRxiPmbhykftQP90Ed5Mk0zcpH/2NLDNFm1tawQHKKkFUAfl5pEFfI2K0by
kJdGvVmTTadR65cVBLLp0D4iQe3+Shc/5QA4oEqaMXL/mPknIwOApypkUs+bW/BRoGoNVxOId2aT
Hwlw1ri5gc61MYqbjzhlbBxiGK6spWnjjDEuvWgDFUHOFg8etenK+FyumY4NUO8frPD1s1a6IRz7
/X2n4hPSWQOyNM1EQ7xtGTBK0e720GnZGIW5fDeSPw6NIMcnxHFsr60NaTdV3rAgsbM0+w7D6+rF
PWljqITvB41+2fmgVvqo5ukq5NQuNNwzEs+gyF/yznw2U/1YlpSwoh3LD8jiOWhIGkBbsBOIomaD
Arr2s4VQNNAvhqut/A+erQZ4P0iNLkrzMLZJwdAPHIN81K0/LLF/n/eAvfK2U+hPUhU+INhIYjc6
iuvF4g2krIHIKNxzSfmHxZUvNAHqDn5eHELHs0O/6FWR5CorA5DsLZQF+NKw2hS+lfZ2j9tXnnJe
QXfkPKLlv1moWK9JHI0hOrQUp0mxDRbhi1V/AroYzTMK+a8lkvc+XatE2HcxvsDGFc3h3/3vtJwV
TSlVdjVolfIEZHYig13mSNrQo5/DBrlanOs0O+VnBl+Uv8ChZZdKBtXUEpBX0/5sKL41fqwqO50d
bMALQcQny2yLr9lCBjTmds1cnwVenRxjYYz5xA0Ffw9k5wMGLYPO3/S/2n+ijDEymqrGVAYhnRyW
rDBi8gaSz2Mx3x1ruVcROI5bUh8871LyS0uAv5HQwiCmx0niU2TYJaiWRK9Am8QWKXsEt0rVZhCh
Pu6+qd5/X4QYSabp9NhC6afi+zxlM2119ygAK7wv85E54NFJp28mdRjhT7FpLLmhJNV9RUOy9Iaz
l75San5DFU3ZvgpbhOXcEp9KTIvtLr6ylgwSLVmuERqIzc+ibO5ul/TuBX8YKY6CycBT8DOZAU6R
CLqd5/jbxsJGkd30C457MLoH7BB19VAML35oulmYY9L1o9du4bI4LagpQmXlpsH7nQuDAasslJxT
tqC2CUA5UTPub7EcogVV0sroPCrh1U1KsGaq+QmJdrtq4J9ABHMZtWH3az5YeTwux6zk551Ug0yo
1fzmtFXC6h3vBr4g7/OQNYQ8Lu05it0ESdkrxpusbQTxsPQq3mtHm8Bdf/eSQayRN7p9GDpPpRyL
ElwW07kNZgDrdm+wihGfnpgYOyzKe+gGVzs6sCKRIouT2Nteuhr/oGqJInNalArl34ifNdJWtEDQ
2eFk+XwB/DtdqbVEfSnt88C3x7mprunbixaqhjtSd/3dGuJ/7Ia/tTrywffif7brgRtypvA0w5YV
6s/9dG0oXcd4hlL/+D5diRXMiCltNrnMzGl7pn5lyt0pVsZCCBHUS/gte1dvul++Q0L+IS4oociY
ros1HaMbPZCJi0o6hwyXX0X7bqHVGMl8lp1odrwrzDScv/pGO2P04wHR0B6Lo02NMTVHmviOTj5f
fSQDaRnf488t8HtYv7t6iDOeipfFdRm+g/eNG0S7gMK9uxAXbl3sXKT0vxD97sEXxqhiB9jScmif
eylCsTvB2CpqGcrUj+RvdrLQ+1OjO5FBLC4gnbLdefNxauFf90gnOIP4x/uWiXFrVU+9wEQaxuFI
v1c59Cgq0gt+jB0A0mYSWZeRt5I6PNE88gFVO50zFjCm/6/2skiM/YbmkYY2YlQmyonT9KNOFnGs
3gNRrBmznfCHJ/yvmJZdiL/qDEZSzQQbKnPau5fD3K9ndXYA3rSK0X1t/NuqEEQQPvLqP+FHyhH5
kOudcIz4zB2YzIs2jdoBa1VQqIGASumCKsIqlBwpTRWCDmQTipkOjx8ayeJ+QStv0S0/2N40kQP9
buM21niirLL1/I8W9BURRlvQUaJ/yQ9Uwk93dt8o3lSahG7DW9YoNtN/suptitCT8avvEJvxO1M5
aSeAQWwMf2CGuUCI5XVj2C4DGKXudvp66myigJZItKaOni+mZKDLH9SVmG3D2PDICuH2R5uEIlTq
e8ez7VEQcydSdOjIJuxxzNyEsEy8V5sr2v9tsql2aUEv2c4XghmVkMBUwniFoTecsSlOKnPSBEg/
Bz+QJhe/ddDCcXbfe056m1Jj55q24As4N6ziDQ+o6Z6oNjpUOw5gvjDtohzKovpxfQ9oAmn646fS
i5lw2urqpGmjKZlczhf92EgFbDEZNqTkj9k2KwyyYAnirSHpLw6+DWDS8pTB5+msxdsgOz0mEKle
2d3E6Yd+9bkud1gytU+7oP19Y+hDPq+zDW7wzByi6eApT5KM0y+rUOkoc6KOLOfJKSxYQ3MrShat
4kNCcQoMWSud18rvA0jTGszsdq/yCvGiyjdZJj11YficCrNhSfnO/eIhddGVgScNGq+1ygNOrCaE
l+IVfxtdv6XylU/O/24l2xFy6z84yUHnxKdnfVk0yACjgEOiICxiE/aToj1SjPxPZaaY1xbGsJEB
4ItjGR5dYbmi1kywDA1jMrZO+XNBtuZS1yZ2vc38p5idfmjVk30FZQRtQvqCkhS9XzFdGPRXdy8P
oisH97BxzPa1MymXZbF7TMfTncvLf3cAxVeGjM8lSbX1Blre82BSoRMGN/qXSL+RSmoJiq6kv+W2
7H/4b6UKGx10uqxqhcxTt6ictgYWkKju/ULBl2U8yfRZ7N0/aLVV1N3gZzEQd2DGGnLb5szVdWgh
ZZ9lOxRO6GDAGtePVQF93s7ZIavKkOfLx4GcaLcw9k5LGHm3UzttdLWO1G5hi/+C+Px8K4CiwIHG
S6gV0pfK7AnMU0tKNtVdGKcLWJTuZGjnF5ig5fVgFL7+ieqmyP/krL9ApyAdyIgVzEOxMTCrCpCP
lFNaYp7nhOHCD4Og8gT0VGyJbBmhqzniGo70iniAzpDmdftluReqzi5biUXZMn5UKEiygOlcpn2O
x7vFsqwJCqJmSCRRb8vule+UteeG0Gtdto2/dGoAlIvh4gyg9vKh3InsmQbwnTdsOhC3xnPVIPZG
numkFTS+Ziuzu6ZdExh4WtSveovT/1Td1GndNre11RzovlYl6Ml2UGcH9T+pWwQ4Gz/jAsxPcuE2
+p5aUp5ZSbo1hHBqwCT8vKcHEw5PzI8BtgCfjcwxiv974+EHMpGgtAlJmsBh8XJ2QgspHscWjXCM
C/aBVq66LA+Kyf7Gcr61Qry1NfNDRBeZ82DCR+OBKIISKryAvqtXIKjgnzuPXsAn92A83xWC2nuw
IHzEusk2UA/LkOHy75p2VsLVKhzIcMpMVdOPohA0tzLV7013E2UVb1th6RHFXgHHQZGwUiJBLv2U
24xajpkbd2MCLGqg68EpyncKzjX2zWrhTgmTWNrqDs5+eKDs0dFNsg245Hk1L+/2SS080Kj4EaO9
VipDYbbknT8NXzIswYWvZX11Nvk7fIOtinzmZSyUAH/+pQ4nO8kkYfPgwGLCLiOo5gSjMOijPop5
eQLDK78O0/CdVhQgDdlVnilY7XNrEGqAWeqXXigrliGr3bgEEM3NRpmwZ30SUmh3N1fEuwtTHTbR
NrC3JkFFBJd8HTaV13XF//q/9fo+xTx90XqzN0mtNC0ZwtJCzlZxJgkD83hPzeQXCC/O/IFaSXb6
z1UEqpBg4u/ZnbVS/MIvbu2DUCrnOAPpUQE8uzP59Vw6glkzrs3MCDVRt7FC+th398ijeNI+7qsh
3MD4nf6M+Budyd5sAboC3IHQS4xni/0mZBh8mkWGsqh2XazxCdG6cMPg3msfN0GV6Y9yjec+NG8j
8W7EFWkCjzPqGjpbsK9TKP4sjE9SpxoSzdljvVkQnXc9b0TwRN5ZFRhbCniQkuvWfEMBcRe8wbhQ
eHv7SgAz0A6/5QjDfEGI7YptijrhPCApCb+jS6CvhfHSOs7Vfc3I9Sixh0o8zJ/CjLSPjlmWS5aq
QrsDW3kmEonEcCOmc16Z3yUS/n2eT0Z+p4J0p8xI+VEFiWYehpzH2jYdEQWIBIqFzLqS+0K5l21i
w5xw1BBfN6TJxLq4kt4H4owNxEBvcpRK5+lOPfshfiLXNLUC0TdDSKikx6qRxkO9FHsOxHh4jnRC
shniN9FgMt0P853Owo8cpHYRxxb9K1nXV5hyF6Deo7dfM+R4OzdY2MySukdNMADvTYYmBCfOKwkF
y9VRZ5PeJ5RPMXOYmI+Dug+OSXIVh5MlDceEmJekDamLQ2Ub42NK8pl4N8r+egKvlYYB8i6UokRN
0A2EUi6J2b5iSx7saK6nnNbobWhat9+lm7U/ZHz4Qs/4ky9FfC9/6/WS3bwqyMAFrpU6Y4hcSARz
QL/MjHoKK32fhEU3YBPdMtQ7ibQ8cezHIx/SDmwPjyHMh5cJLBLAeAFMiHwU/JngXT25UT8eEIeA
XkM70nKsCqjG8Y6DW/ZqJOgIahWdHyf4NWwOErnGCWWL8MXRFB/2endnJ7T/Epc3TdICKCE7Zvma
pCLwOVzJ9XRQO5VvtGosval6RNjOyVAQvg6nSS63F+bCj863wJPWNGBjjUdAQXxFmxf1GtNHvige
hAiA+YrGD8hK2abfGIOdI97ueHVvSpWNZS1oSqnua1EMyWtcT95HH/2rY/bDl3kVuLhZe/bOnWn5
Lxs6EKQryVHmbOfJsIuckhkkCqbxuO4wg9b0dR+sURLBRJ3BxZEh7ewc9oLc8QfPcBq1gzvbvCyf
JrH34ZXa6EfIIgW0I3XjDeIdUmJxoc9yiinJ91lFp/2/kr/j6GLk4zLcnzCw8dlgvxsaRSJ/gK6O
X/VXImWFGPHwJkp81xk29o8PLpUyGB3CaqfHdb/kfRhmCeJP2eK0gMKvkyTBrWxGagoLVQ1mnTNT
no8Y55mqUzZxWd/ITMT4vq/wOG+yPHlIFHEsdBJ/AoB2ES9VXt5cC3TKSNw8OIDOoYjh5Xr26mYu
6tkZPmu8yoRhJ4YbGIV43QXnJ17fj8pZ16oV//yLbcfPYSOJ0gsjdsqQw69Dn1VxIZDmTSCyVhWv
SsIZNEy3EWMhHGrHT7uhG4m8Fxin7OMioN9g88Y7iU6h7kQ7Eq/euzsA1wgE1uyT8GVHq7sbYO0d
RkPdAETQNCotvNkUDhmqQLanH8aVAGbZRjSytfeNj50TpTj+9oFMJtbhN+cSHR+5FKh9RE5M0Ip9
yQ1dX0NVtL1lZpX65B7F3pCg5auFgW8gjmpEugv85vS4k264H6TuSzWJ5UnCXqW+bKVg7l3KP0rd
rlBxcu43Vm56PDlPzaCJ2wnuk/B2Q73njlKRspZIr9mA9XdPfyRKsR6nL+fEubbPJrP1+0HYm3hR
yQhTrnmBJSaklBCqx1ogXyBd2prDOfQQbjts2rzy96gsbXTzLT1giHe/6MD+jFEF/+n/woFOHyrk
do4DK0CYJW5xTJeDzp9uVSyVzvguYS1ID3ot4g3vfv+vRyu0U5AET5Ai2ykMspY6BAxKiRDjSEuL
tFpUMApviJbrTA2pW2T4uOHxQBbb+SzavEW7XJkA+6woiVKjb76aWo7g83FQiFyW+5CzVn4dUqVZ
J+HmY9h3XZ40/zAbezA96IZQO+OcU++NhEMmS78Bud9mhdBD8Cs79VBgHPqegqXYAmUeW5TPphSH
ZCDKo+uu/XrBSw2MLdFg04S5ia5UBoWcdRSUNIpTcHvbUevEv8QJhaN20nKXpTamppJHi83NY5Ph
DqgAcgyGJ6AZI6INrVwIZE7yDkVXvJy6YLb6JCZ19Ot2Klz5sQg9Y+y8uRyo4cKGjXE9NLtiMmtB
sw3jD6Y6X3NyxxvT4xu+zi6dJqHIK2H6QF0sX9JDcWqGuMsDN8VR/soappHrsOSIYbbWLA7h7YLA
dXxHx+PNKkQfG0Gted7AszbwXW2TaoC8ag==
`protect end_protected
