-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
uGwM2+dGVEnZmNOAvMgaczhyeriKipPHIRuJo2eAqnfCsX8fc0vIN/o5A8CG2KPF3I3HpqxIRvEk
QEBDUBeRv9db0896OIXrkiuDZ1qWUb0eEnG5JDahOCvwRbDZObRnbV2HKBhRShNPuVai/sgWD4/X
MTo+Avr57q6bZLT1ZkFQAJjKy2ypgqx37D6ouqBHwReYSfFkYiViGLrL2bxH1/TmxPmayz5V8OOU
zEqBZQv1TfMwym6m1e+oWiwb5fs8w/llV68/YBdDH9RB7018iGlkChnbJeLc4qZhVVuGixnMH+io
WA4LNfrCVPTSOmQ0/LrCM9fAlTZydLiuh6klAg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6224)
`protect data_block
/dTyD/IocaBnMPaogh7lF7GwpunU6M5ObXrtROfVYaqGGXj8njAkokM5ZhTP33tN+J53d8TP2abJ
9V5aNnEAPnZww9pYzH95rzunBTF3AJXN1vVNDw4n+W7/rs3TdvFZQk2HSGWGrw3UlbRiGHzoJokb
oAVGMYGtmgJICDjovOeX1pkQgGxay6dllprGy0st4+Rr9CkALh33I+zYpxgJDJRAZWgbnC2bfVCY
GpVuKljSzwMYbs9zrvOcMAvoygrNyk6CbQWOPiQd4v5/sA+GNxNpyvmIu33kazJvYFJv6dDMwzzY
xSGESbPHiC/wR6O+KcMwv5gEAD/ge4VBtVBMlp1i3fungSlA+7AJqhdLAkNmw3GuRWfSCAtPDJ7e
Dw2t68vXWXMeBMQ3Sj87ARNRVGJFyCpGHxg8vHnd8edooZFaZl4UqLdf13YZQxWumr4kI3CvlnOM
eiX8vY2x1n8UAEg/1zqohBlSucBLwzkR+ip1HqGZtcg/VOrCtFykdXWHUr4wpAV9si/ZsH/w5+zS
wEfQK7YxtNiGpjp9w0aTew6kZ1GHBwdBv+Qk/6NJCjTch5QIYAWYA+XETcl/fOBAgMnQsUYBzZ4w
p31WwN1F8nrPKXTirPOFsdwZVH+X9RENahx1zxeQGrBQ8m0XDWqR8qSm8xQ2o5NzhHiyBZbNbqn2
6m/WmeTyMShmMPCTqugrF/6k4+0N2mHWTl9KcjVa/vRwlbOv7URtlD9fmg01uKGO6TQXg74WR99t
qtMQFTqeIjtNUY7sjzfVMhJ3zY+ZJcZNLSfMIRxo1U/eYGV2bZllhWj3T/k23dK7lgD10p8hHLMc
ZFqKXajkRXi66hL+5W6Qsq+Wojodt9pAPqtq95SfxhDWM/wWUjBTFecIIjPfHp7Omv9AjfNJs8NR
cTSDfAwyWEumoKFohO3xwWxI8psls8pRf5CJWeneHkEFfYulcA1ZwolWc3RcFNufbqBzIrZEaXSK
19ArEQnBG4K2LeAmVPr/pZibODchDjAEztBp6wKgD/lbPBQ95hF+9Iv56v99oPpBuA92qT23M53X
haQDagxP3FNrZH/2mqDwbbkeJfztS4CuywojSwpNiEGntiq4m0zi5qOX4V/qxm0suGw5KVbUcTlp
izpyaWhJGcCOT7FiiaSVE7JlPR8k7+xTSoC4bUtXqJmlc/chZJTJmLxxLovXjUhSVHPs7BuGyGPe
ndjGls88pasH/iy0jvLa4BoH70ooQGuBj+Y90/gV509AJnbccH9KiJcbm6hWCJlWP0TksH13nWux
/24XjUVM9P7RBWRxqn0QHNQ03HNN7WB8ImzAGIkx3E9jtL8NnZhfEZcxzDirYVoFJEPsh8Z7aVdB
298V8AEHv/XHKzVhlkI65RS8xLOjsOcxLhtLQ2MTNcDXjpJGk7boB8A1ZdaNil/UfFRLOEUBkH5s
3hv+UYTwQ7x/Z18v9JFHApUQphoW+0A9VC5/rp+uKazwSYV61TL3PKdekpzeQPee+wzxCHIc3VtA
QAzS3MKlfxBnsX/7wrDwXCmrc4s8Dpd2vjyGbZKdm3g7sI2K3gYAkSuVJdd233j2I+E14RCfBlPm
1KBfjTllsO91ng6VqJ94AFCeQPIMdishL0Lshil+QOH3dMO4P3YIooU3x5poMOQlTHA0bHT9z8dN
aobgXCS+TC5KLwQx2ic30446Td0uG4AgiLtmGdcA38YqZz9w4qhN+QemLN7iQjpYdLnbooeUaQ2I
NDN2AU0HtqoS+aoHWZqFzOB3XE+yZ1FSscSCL/z40Qa5XL8X6XEsWPAqHB7yw5jLwpmJg2dzy+PZ
d0xEdONSamlnl1fFoKgRRkxylsK+diowo7EZy2lFTx8eJ8p50zNSLz6kzNFPGe9hSmTTIxiyWTrr
EdK/ApEovqdQ4UZFtnFkR62/cdn7YYYgtIP7q1qh8Z/jiu0JqNLpsGWarcYex73L0LeqM4xcvdM5
20hKM3+r7xZZW3MS6tHrTKyIES15NET8sXBayRKM+RL4IsWpnFkA4g2oGJZot/bUowQWHmKW7OgI
82TGXwGPgo6J/QFf8ITbgKTXPXvESbkTYJeAIh4LVGE4PcJNcSxnuqSwYkUTc/zx/FxyIKMQ2b2Y
8XhGpbOMjY5CVmEb4pGYoYZhRWbNnaJ82eHPNa9FuVNSaHpBlSUUQdx8fUcOCpF7NeAj/4ZLiJoO
HRlB3/Ex0rMgbcRo5BKC/1WDrCX/TbxTE6xtU+xmB85MqXezKnyENTwa9WeFfe4QCl/Po75nA8ry
1W3fmWt4xAtz8VbTUsjQYFi0uga5qOdvjwsC9lREFWn1+6T+Q4b5lvIT0aVuv5ohRxTuVJ6z0Taw
/Y+2pazjSsAxvUOHDzqDKYIRN0cdnnyDMgBqxzKCqAmEHvbZrI5jsoCp90Rx8BnHUgWwAHxJFOpd
v+YLbSnAJuHDATJAs7nHtP9PsMh+A0NDy6EpGo9ZWq1WpTaiL5x1CXqh/rWLvUTU7nd8xLMhB3W+
CoTHM195prPb4Mej9T0UxDsaxml4bM93O/IhZK34llrrk5Gq+9fF5KAOIjiG62kzpr9AfZXnHCki
KVvVtW9yBcJxv6nDCu0LDOoeVu4f1moNHnBNczjD7CtD6+gd+Z1qgjrl1FJ41dIHfXVw4v5jonfs
ASoaNcwGxzcCMdRpFas9wg8DyXQj+CBHGuoaIy9CvtEWqSMY9w9D0jx2hLn6KW7zCx4ok3ytWHPi
k74PYmMovHvKafdtqA7ZB1TYyvbcCn4OpK4kGNFTXQ7UyeMTJUnSrHg+sMVKvNXBdlb/3MDpGEGI
Gu2aN1ml08S+e+OWhgxgjTBaU3VcF2K2MoGZwtnCwozXlEzYpEdx8/l2Fi2+5/VeLcr7+X3q6lSg
ZsvOlDaDcsqUZ9D6GruOggJtzXXmemky4YzAPZ5n3Aci6uu2mb7tXuYGrtrFdPewbpwYibr9XnEj
aJsIiXPkTABZeI8LBaYqh1hM2OLGkHP8r7WhbsrWbkcfGWExyZAXD3oePmj4bmpNr+3sSg9/xXPi
6jOXRoVHCdQ0tyZgyzv6L+R3mGm84dGUhsmVNeLmBuqruB10iOfBF985zi/N7T/6w2A4ZfMbGmZn
gjjjB/GWyidffaLh5FuIlRy/WY/XsjpTmuICCjHAu1DZSJqPEqfMAf9OP9Fy3dwN4rrPPYwCEIav
QnNXk6SPM5MkGcPrhYXBH+RcJhehqfabloftUNhYvu9rv3xEA5u9w57lKhei7KVQlShZ0MVJAhmq
u1rWwxdpbkCJnB8Vkhfmjd73befPMd+6pBfQJZH0h5cLgKxkJm33Cu6h0EdtsqmMYE+Ca0PONOwD
8KIwni/eDNl2CUYXpLlJbsZGsAZ9cp8CtLSKmwgcm9HCWwbCFrrYcJ2nDExEDpPjeBirF/fU9gY1
D0o6L3A4g+XKkzQlFwq/x9gR3Z6Elce6Nsya+feeBV8tcHz+oRRAPP8SXu0FF2g0WhVNwqsxwiMl
d0ie2VwNrn9ayU2YeChIC6a6hSfasBghoSesNhzDkaA0schvc1jrr/M4aY1VfZZDIKld8PesxhnR
8gNogy36Yil7QXmOQoWS++VcN4ZCUT6jvcs5RhgyEhHBoVYUEUgMCgOFR/0eWvtGYSONiJTJ3pKu
qANALovfWw9JEEBHDwqWbSu0jZpNbdZ/IlLNtdhYALdoEyroCvj5H7jZgYJH5tDuwBWttDXakuX2
MfepKZ7G2ZdGU6wMykm/8n6FfpJV7lYNIOGpFeDwC6mT+dfGYs6PlgizZj70preETHo3g4BW/835
ZNFi/KOBobDa91E8pbz0o+XRDyxgcnvoFX2rOATncF36HusubO988z+OWeuPUlqZtLO9NbXBi5XU
+GoVFtsMaNKb8A3vYEd21kZseVzb1oNKHF8v/NcA4T2+iPBbOqSa65fZeUj4MH6K0v3Cb0vJMvQd
DU5ghbGIopaOEOcM7+LAFwQS0bKWyNUaCUzw77kVaHGFyRbTuHkq1Fe29SCArZ74vPUFJ0zW0NNR
5PovQO2JGEc74lGKDwfdl34tJDGbvVOnhzEcxu9l19khKOUEUIGgPzeE5H2RuelnZlGWqDTOoJZS
Ied1CFHptRB2+P1uwjTguZTr3Uxyrb0ym2oRHkV2msH0TLzWIp4zelvKaY8huNg+VDYh0D1SrX10
D3PGFeLIViIUfahEp7DOgWvAuj1Pxew5w/AtKJ/4loWpwFm8cA7Wn2RLhoeUExo7Kp2JzoCodvIM
jw62eTNrvzt6/8hGspwAu3rKhlg83wpbsXvUSjVGex64GQHJtV66tR4Mse8c6sutD81tQmzZ68P7
6jnkzKiKFCjjloUUnWRe7j+/dxM7NeXTRuL0IkvxhF9S024snnx1oK5LZfjS4hhUn8PpNV8swKrt
qPrDicnkgJPOZEuTtSzeQqXKga+DPeVbJQjt1mkIKkSRlAT6TPyA0C9JUJ2+pWy/Pwsx1YiCXK3A
yGuIdUxbZ17W2h06P0mylORl5Lkp6RmnBSTANrPAIMT6CVWzR0a0nv0xY7nudmNnzy2VMbNBT7AJ
21uJPNOT8KvCDV7j46+nZ00LkHKjjxJeY/n4SbTusIoDXPwtv7OvG85taiKfgXaaHIBE+r3Y2Pxj
Tyh4I5ny5cI5myg2xNHavjUHx/t4QYU+KXuAdXrdyewuaIroTcn6niY95Znk4reIfatPNuKZDurI
wXuYmEtjPhRaeXdrWh0URODCLgqMzklzEbV9z7htLVVoSRYB63OlYgLZAzHx0DNahQmxyI/6FfLi
hxBF9PjAmaR5Ff/P1eBmEn6BKlmcS13qJsIk6B/R00C3pxkFwyedu/CKVexJZ5RHpJyLYyA6+iOa
ygvWkhc/mk44yY04T1NEpmWfjd3CBv57E03YbE6MsaU/BHyFmwh6cHCHtDQF9FAryXdHXk6zRpIe
2koDot6zgrsWNF0aBFlCqHIqO5jg2+zzHjBa1YfqXvBNxivaCwt7VUu8lFyy96r3GLe98dI2TYgi
H966yQji2BkuF7KJOlRmVyuA/Tl4+/WyWUXbAfcbMKDoQHFgWD+8sYy8iE/41ZdIVmTCYXOVGphB
mf76yyXkBXWboDh/pQVd5xhQWhkaddjf+xaXZx6VzFqKOUn/5a+Gto5eemvaEGjcc3H7KIvkejTV
iHq98FA7E59Ea4uUqsEkE+RSgl2IGZA7IHQZPbS7rq9jPzDla1vMN//VYmCOuvspVynU9tDlfd+8
PAYc4XevvZWuanjvpeBUtDiIHBF5Iqg5NJJWAxP7jtGrk4WVHK/+fmSCssouHL2GZdGS2qUQQp86
97XkWXTeps9/fjvVhOBvz4Vzs+LGMEg5m2BJ6i/e9iX4VFnu1dywiP86RcUw4AEpJKrsrL0flKpl
UM8UnqpkiJE2HsMokBYUpcpjBCT3GjKz5LVBWDFYCcNlTOy86aUv5bAb3i8YWH8xLegiJLomo7Ag
DGw0++NpTwIjh6WFd1sJbHxtRzDKWglU9nO1YTCqagDhqlwpnuLZa4asvarZNU6iY8LjjVz3EnkZ
IeDIzjXTJHR6biyRBGEPo7Za3PBO6wLuVhBIQ+rRjGln9oA9PKSBlhjEUzXvEF2NORPF3eDQiCiX
jrTl62mCeRzaQ2LctdQhqHLArfnuRT1oDpbTscMkTc76W+qVDE3FpwIf5qmGybNjeLKfUA2LEj30
mYtMQ7BuptIHhxbay5WCM2Nhm5OPPT54zAC3KXON5pofIpCnlch5TjuWp/sJISt5zevjLGEBkxw4
Ve5N50p7wMld7fMkUos76zHBc4LuXd8+wid7JBmz+Zrs6INP8STl5WyHVxpWO3cG+TLJhbmEf1qZ
G+4PKdTnHJBjeT98zU1+JC8ZYmL39pBA81WF4C4GPw98uM4dypnRGD+BjiLCyzRldyXCB8VlHZZX
kY5c1OXRI+orOUvKEk+WrNBKUUnG0VyxnDYDmL2w7rQlrpVARYYZ/ekPdtIR2wug7Wp/WAYoGnvJ
/Bt1Bm+nbzjdp8Y/9GVD4dE5wzaEjdFJdvZLJDEvv43FoJH68h0033uyl2CXa6d7rodOm4Tkt2Ix
c+ahNarlaOZRnkj1a/ZIFxYt28Dp+CmrItTjlHT+tPV8wSmpjIp7pnP+nOJR51ItRRIXdvVrq+u4
FQD22hIAgMx3W5RQyKrduhaWfOPl21zKFpbpfPpBK728Aipl/157S15IamQU9rG9E+ULOGGpj2sa
GwpewNFzXjYR2lsR30kk2PnvwnwDXLZyNaaQT3/TIXJEPn1rcDLcGBtZxXCLLh/gQAFD8qOi4glo
0MQmxPUnU6qT62SaaoRzAUOkdDjFHWeYpVjtgQvYR+l9ufTW2D/rfBi0IbQ4FXeIq1uN8RHqFU5Z
2xMk1GMMlMH+yn/h1U9m31d834zwXiPzij41fifiu34IqfaVlBT/Di4S1GVpKYu0Wv25tp1nRw03
iB/V0+GdQ6EzUy7BMRzYo20wcsuU7BFkTGUrT5Jk20vlky71PayEkfIw5YQHsH0c5brIUoqH+l9L
D7am7py/ZTMsOo74CxRGJcg5uGztVnnrOCjFVnHwJFYdIudt/c8PKy7+GFMHpAWXKXWhgtttLPMv
1rEaxftZvuHuTwHoTOr/O6LjSg9a/k8hNic4bNxzQ1TLef3l5z92xUG8ew1LUhpZ2KCS0iccrY7Z
RC5zTz71H6oQPq++B7tVU0YXyOqSfSZN5voPCRja6EGKCT4z+PgHdtKsIrvTYXQlye5qwxLdNwMS
nIgh85P2KoQZ8ci5sqF12wQtpJZpyxcKTZFV5929V8SvaFqIBFaMyTZv0rrMJEFSrY+Tm1UZrzn8
rZuWZ2fMCDbDhlPsT3HpWOUA15UOR1joIy8N+ivH0nRcsQFLvSQWoL9k0y94xlDPzKS5mzJwbhO3
fdI3Uqv++0s976CtjZsKzkW0WWOChfYGkxYTELxiERxqkRvnU1sqMsLN/d8LSFCjoJhOsZOApZ9R
SW6VVk6OfXYKladteds/STjo5wqCvjTiSjhDAQE1fq+xyPfIHBmwLLKeToZAZH/TwU20tsxTS8mN
M48yR0wL1P8hsM7cbMwamANhw3SYiQznqYPr40mm/b+ya/281fbuGsqdTZRAtfr4nbxEI2KFkDP7
iqedc3OOl8kJFHPSUUcCGU3TJQCGoprdOnb/GB30xnFmVpgGnHVK+BlRHhjghmfWwW4TuCJs6gOv
4g9IMFQGaxezwiBH3ZxTkPfUM5ZeG9eHbFxg+UhYGMhF5dJhuEMcPyn5l5JebSYHGBG54C2F6T0T
8CE4bVXhcG6Szq9QdhRgpnaDu3me3i/iPXvkLvH3aC09DQs6ZXhf2/xbjOH51dHILO1m/M3MCxBX
cEKIvy0BPYylOCdGP3EeBv/ZeAYCk4qrU64Kc7dd7WNZU0oSFmXz3c8jxYFV1K+hkuR19UKaGL3c
N7NiAPzJVZTGUeB1RN5q9lhdLgLsY87ztW9mAT82fS/c/yj0zTd2JLprCjeK8W6tdpHPxdnLyPB/
V/LUDTPFDxohuO09zfcKbKL1WzbnrN9u2zi2Dh9Y/nl+zGPfidbHgfXMh7KBDPcU5pWv8eZp7y0u
jCIGUZTUb6kqMCBPuVPP8OM6hsKcpH/Byku3GLu5zqEQP3MS5K2sh03gdIAZ0xlumVBOG0iFMDoO
gz7+R78TwPZRyXuzgjq0VgZjLWMeeFdAJf/cCDwgMki3vCCLN6ibcAcK8KedtfLWi/q0inTcyMtH
u+m8gWSP59/N+4PH7fDpOK59uh94dqvKDMIofbXRrX3wg9ZOkZCHUzTSlHxri9pRJjEHafQL6gmE
Imfk93xmdY07HmIxIYE5GL8Txk0k/zsw1PyxLiGItUtdMeQ2GXpv0SVr7hvUknK4Ijn4jgKCG3nC
LyHCXJWpGzSHF9HAUWXbtsKMt2Xiinfb2fvAZAQmYi2uicSLOKMcer7Tf8XjnPJKU8zwjQDf+eBF
Tn2bbthf60w9h52Pt2CY6ToJOAgb5gj8bVC9LGhoyP/RKNWVnKCXgvZzAs5GY5Lv2LxSRDdr3KBJ
zmYVOSdRycnPK03MmnzaAHMPDsf2Sv45OQ9ihcebIz4s3v55tJzVsVuGDztEjYGM5aSF3Jp1W64Z
tsl+bhSb8s8X+W8CtA6uvcv4C1O58Sv+Y/1ZSiOpRmxYWNpbUK1An7Ms0D8FJQFX5Ni/8rWq2mu9
klkBBxRbiuzOg1/gELKlOjPEsgWBZgIB5BHQruqzmOdVLJ1h4BJX1ajwh9dnwIE3v87uxbWuIuYE
dC5i7SnWbXHDANo=
`protect end_protected
