-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
cYVArNkJ/HeDHxQNgHregHbxFG3RjuA3eZTuBKHpKhNUruP5bSEJ2C6RhV1hC2NgYW5JMQBsA48T
3A6cVL5CxYbk60sT4YKFxo7VF/vqlfKwfj/JNRVHf6OsurVUpTVJgQ/FXzhIo4mnK0Tj5tSUtfIF
lys/b48Ng27fM/4Hmq5sAEOj45JV9V1cdRhhy2QMHz0UoASLvMp8Vhj88uxcAiy8mQMhGxTeOoOb
vnbqQ8jUZZFQZfCgsLRMRbDgmLRdQXi5JpfhRNEy9RtSrdrMrxaiPQiQTShHYz/BbDoKngsWyFje
g1mlgsmVE9xw/j3PqSVh27dbj5gABpwMwEKgdg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3328)
`protect data_block
ALrAGIX/SXpuBEkb6QqHKL9cQdmxVpiLweaNgEcIAU7EA2q8R8F6TZaMfjxfhxCxpfzPLxYUBffE
qELGSw0jMqb+g9v/F0yC91WrOS33Suul21obq4ViIkQpr2mIw/za/kF9H8lu7dmigK0RfDheM5Xm
Q/oUZSDXhKDOv2uUuN7roQ4HTOdjBwxbNg4kCqBSxA9Qz0yK/c95HiGx7SMjvBiU7RrsvhtpXhWk
dIKTKBBTR4/JKWMURpugPmrHk64Z6pd+F2sw6q+QhtVEPIg7/W1bT6eKOJv+zoarc0bgQ7Swn+Il
lGj1+d6+gwrv9qXrbp7n7xjLVl8OS3mzm00XhlmYXcaHmi1biXd80zCTJQTTDIjMxVaoGaGaYa6s
v7aVRiTBzhMdBCHfDgsGhIRbAG6ScUfRblcbWxSxAKBFYwfoYoRUQjrn+YGfX8cOeGg6HhG7EZSp
yVQvr1IvEc7dFhfNxsfWGoR3vis+ruTInF8Pl+S0s/mz+AxHUzSlWJ5I0BNHbFg6FFl/zlGuKrXp
gMFyxo43bOW0LCs0nKq9ISFhaRTV+xu8J7nuzowbCmwlwtgCbneYjgqgFNHHZTUS9Y+MmAshIckn
/UtZsotLzt6hvarUg0EOSF9XJ9lHemQFURzkRMFDrB7k3RqX8r6gJauque1ZAuYbttAzxMjSSDpV
DKhlARlSyPUq7Bz/iatenknwIYlt9an0pHQVf5Hl0SYIKoBsfunJJBlpdmHw5WBaG3lOwPzlKFsU
pI8IqPn9iB2nGc7A8v/ie8YSRck6l7X/lAme7wrdHailWojgsezqCTo/Gv0IP0bunLIyPOTpQWGC
cVyhn1layUS6uK/YNsz/1rQyR43CsE2I+W40ePQlWLJaQxIIxwAEakB9nvgSa3p1ezp7a24JHzdz
mePYJQGJY62hxrpz9acAD4OovY3SrMUmmjVodQLrAi0UK6out2BwRS6BAEviTva5NBiU4X1zwdPJ
rA4KHGJrfMlYA889e0JhXCHxZdJQyNmS0hxHaAc+DVbawcTOxUzDaEj2stiMTlRGqpYJsmf3fIjA
Do2S3ULsEkHew+aU/yMAjQSj+vPezkgB4mRdT9aYQwQ1FyEgp/9hgMFiKWwefaKLjQQ5WVmGi8B0
hDlNJwKYbnivk9v9Fm8KceFYmF8Y3Y1kkglL9oakjztco1gDgUhSY4ajAConVpDCAzQW5Be4thVG
+L1hk53yXSJ0hDUR7HYRs01Vw4NS8tXQ+X0DQjv0ZlmIHUyPfO8f0O94jaxWTq6C0reZQed03oFJ
KugmXJHFqaLaoBTX7QR7zg9znSlUqC9dirNuLSogmMk6dLkG96FWRf8Dp7uAYAchVoLG0EdgWdjv
ddRxMdv2zBlpN50xLD8yDnuNmbqL8PwFKc7dFFSS/l5OHYKwgWiWH7AAYG3TSauvE7ow0cjc3gV3
kC5xdVYgJIPB60SABYiJyXOp9NXrbHjipWWamZBwW6K1eaM7PryBItYfjJOXAmn9PM0laqJYT3mg
GbdGD9Gvdj0x1MWM355d6Oa5XVladtzSipQemO+syz3qudbeKBLuWjuuLVmfw6SIeKFvag19Z1of
ctCDtVEMOBSG9kSAnSDSDXAzc6TK/Mz/bpYaGaKOmOEd/R2NyTSC02PnkM79typqNneaC3m0xy8y
4IN9mv0immHDj2Euz2QUPYByPJOh82u/B5Jypg3m0XYQg4U1r6shC8a6L4Ob1CDvTlCjzfcO3Nat
LkmWuEu3Sn6TNqrWmCPhPj6XVqE0Y9YaLIECEXd4SDJjrna0mgbZ3en9okWkaaJ6JvI+J/PgLvu6
Wy3Hd0NQrtoFywvIygLBKHRguwA8nV9qTFXXa7yzDUPh7TKA7mjnmw4N6O8kIoTdAkfIVqDwqDOQ
L1h9E0ICShdWBOgUO+koUNkoIoA3FpEojwFALQt1Nwy1EhTA5JMjBgSIonq9H4CdF7bhXWrOpCkR
q6ZLCRb5PE0/ZX5EWVVqHOU6IdfD7FUj1//TwrVv2Ts0cBYADX6/tQvkn2QmmS7F5Icind+R14NW
Hrx9/KCTowE1Xkj2HZkD7voJAkZjwHKSARJZxGzXvkARRtOTvYr0TD8lkKuNOrrMhIAp7yn3+3zX
N2M3ybZL30m96xdhscQ1dbQu2sXHeHLkuB0YCSWGOTf3vo5MbsjRH5LEjTr4y/b7xJqUr6LG9uuL
IfRDB3gk/o/3ucdLFDzDddRadg1xL2yexr6tsrb7qQ6dAmiLpzQ9HKWRiPKs+O1+kH2TPw0Jsyix
PN8srSBphEX9KoaAkCXNFOGLnV1Q9wAc6+qWqTkpLHqCYdE8BJSSW2zpZO4O25T8z4ETdM8rb7TM
KXo7rwP0a4sscM5eu9MZfnUN/cH1lPfS3W5K/up5H8l7koDSYRhXqUIDQ11FSdcl/KQ8fES7wHaO
3TlKCi6efBos3npuh0BXi3nYU9C8jmrZ3CiutRadHC7Cf8A8Rqx3+mxwhtz59NfLZ1fpVWRJTlU8
uoC/H+4TeNZZFaORmMIxxTYlVd6r7akUBrQJDBpvV7x1KhYyRcOxPsWhmzggDiqguIgbfPUcQ6fS
6rJwhWF62poxB0/6MjOQd7cx90tVYVS9hoNo1/EaaqpchLB6ldKaOCXxaTSdKYSKxzgZu3mkBbOB
joNIm5MKPDFFls/qCeKbJu918TYiDbwp/yp6oEEpkB+D0nyMhBWHepmVPiKLzQjK3DqLY9jhMOnc
M73UZv23UHyzG5eQmGZVtL9cuoLHDVWMgroYkTzBPDk/Qz0ugWCYkdWWMacQsG1tNefgLhh9lVuV
Kpf830gAoNP0fdr35EeYS7374zmJ0yDGxWFAxvgIp5xRlgy/IvqkrUTFc585s/BHCVqxEhFVVs2m
KEf4KSU0YdeOLf+3bBhL7OMeoJNlGUm42+4S5foIEBwVqxaonuvwhFvB2IKrRNKwSVV5oMbHYwyA
n/vKIqKID294TSI5ZLNNUX7IJwVJyBTDTv/GyYjXaDOuQNPLMQQ/0AKqM97LZGMTprc9JVGhPvGb
iR/HEg4cv8M+IeamInvTLW8ox6ZUrwqDq17tJxvJmP8OENvpG05Xc6RhQ1R37HaiWzVKOMLkrkRj
XTBSqzMa409dm9H6Vkv4UicjckoIFOyffIc5Zronv/P6C9bsghDgMLtHUbQvP9goFSz3710vv1A6
dbXC8Ogr9dFL5+99NCS6ELYwsClvFIrW4XgykRLorMopfcLynWiQIKychw/SbYxVFNWVem/e4zUE
coVciOjw/9uDQtcqX0DCQELRHFy1wmfNXK2B6A3XEPTfOlxDqvWCdHJQzXN8dXHqxachtk1zAJXr
7Dlsm2DZWGMlfPi2idYJLRtvM4S33agJxL5g8hbiW9xomWPBNKlECEYM7KeHHY6QsmN6CHCRVr3o
In5yCR6XtY0LobEkZSzjFzu1Gj8arbw23uevwjmTRRFRANp9pykXFvPv1MVEVbX1JOxM3S2N91Pr
jZJeO11iGJ4Pg/Dk7RQq+6m2PT235uFG3HyVT5xir74BEF7cqZO+IPbKkXtla6cgBiP90js2fzw7
3hI/m+s+tL/0FxDOO6mNc/hcUGuCSFNE39czzuiXHbLjoEj6cox8dVFSzgnMqKAcFI6zq64OxFPX
KG333zMAHwoGcw+yCjrbc6LZGnDHuclC4kqqbKoyk8tTPg0JwzzilOOEidHisi050GGaROiUgyUs
qzGY8RUN6nZJdI+Y6uS9RzkyjBX66L32GwyToSDVXX233HItqL2aO10USa+UJ0fISEegECeesCl7
pBGPH9cbMPkwmWKViIPTPtjqDCMYgKbj5gq/L8zXeO9WAKdumtDCAEIkmyhYyMp6CTlR6CtrFgKc
78hlvr/DDobPfW0KX8N9hVeUY1Dsw1HtmpXPYt+JDzR7tYZ8G+YgAYRTpqETv1o5Ts4yaFaysrMN
AUHET3fknHSP1mxtmAppDvdbEMJlL6ZvcZLUZu28W1ukwElDFq/cgl+GEtLI3tstgYX6adjttqDZ
Ha/XhfvuiClMJpAwgOP8Oq3C5EO4FyVfeMVHTh3ZxrdExvxt4Q0ouCUUdtGHHDUA/tnC67PzSErR
S+sNCFxnm4BCXiFME/dDE03K8X01/EnAQWsGw9Y7A7+UHagce1KKBTHDPL6PaPzXJDPv+fIrewi6
m15zZGHqIFBMar5FiHqduOVgNiWiXXnxIJAd1srJ9p7PNDJBVdVoakoNjFOnptL94Ehlez5+ZkbP
njRLPhHbmEJxl0A+WXUIKFiyJHcqpibA8GA/l7bICUF35DdIao1i4CkeYAmfqA/JDu4MWxtXtyBn
3IcZbT41Cvonwsbq9RKaOhFhvF76TIW57r2qfT4RPPw3Xsiex6/x8SukmeR9cax8qAwTMRUcpkB+
a8OSduzpmAss0RgdUPWgGFZIh6p8WQ==
`protect end_protected
