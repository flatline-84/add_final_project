-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
QiZgjWA2JmXdXC+RCnanuosjA0zqf5mx5nfQ43o+mC0CJEegQCsnmvSp07tOpzCzQGde+MzseqdE
Y0rP9dhT98H8PBXNzfxlmbctRonnbXXjDNohc527ut0O+9afzUJ94nYqHwKYNhKUDjmXtQGD9yOS
e0czozigEtNO0X8xNsQo1tO1k9sHXsGLf6Rfw4nJLcoWipMB7TsVZzwzdFqIZ7e1RCwWTJ3N8Vs0
5mQTgIDmAB8xEEfrPr4QQRWNccyMgBI4BzvBYXxo1L9iT+hQYSALz+hows7efJ2jX19WIH0iqB+y
V6zBgYdHRCmLHz3yL3jd1VpGEvPIOZZ7b9uiPg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1728)
`protect data_block
r6bOFqY2YdhIN/SaypqKTLuI6D1jzLBVq/bddHarQ0HSQ6dlDlqe4LsNzBvTPFL/Sij3OwaCLoV+
sb5RdTZQ4uzUr/w6fYvG+PknCIdlNm9IN5fB8DbafWnO+gsw69Y3H4tl88nYhyM31yZ/L22k7zF9
mkLtQu0W4q6m+Hz5viT2iKC2rCRbqrL3ZeTu6iBrvvySr+MAL+t1uj269IWzMDZYXgFsmiHAKfnN
BJY5Rdup0+3yrVDJwx4sncCL30/LBuxwsV95W1m0dYtWLagDmpO1CpTMzvWOTab03oYSbgw8JeuD
dy+0iiP+POZAPtsBsjGNfN0Ukb2xjV+BGOlTvj/ekrKJj72lMnpQhjU2CXfxBXpCY9PYzIDDL5eW
9QWwUleaZtOuMk6/wj4qk1hp/W9IxYDncPimCr5cUYvjAQ2BxFGGSQ4txNPp4tfEYNE9LIaHdoqi
HpzM+xmCayHD3kPHn+4/1V0FOZnKNZisZQ+ikXDtSTG8r4x1h4M2mgibqzXFAzFJrZs7bkcbBdSe
ruU7cHAV14sVL5tJCmxo/D6TkkT7bO/5nxZ6PId6voa/oiRsi1rg47M2iIghoxUpBE1x7jQ94WjZ
MuHzoTMwWD4uTJz8dXM14h8Uf5Rnl4vGvPyfV9mwAnPgfZmhf2rLKsAf7vMGvmBpEjf4rv98Hodf
/QACOzRgIFT3MsBjnvYzzK1v7r/JX5v7hWRxGVZvGMFQqPtaMyUvxCyz6FpTJP2c6mvqDaoQoGzk
oHd53CrrOqEU6kPMUoqofOmorbC7XIntVcl3GUPMhm4LEjUbQSii4eKmzH/0pLsmPBL9yHYDaBNf
bsR3P0Jw1WEHvU9fsuhVPjj8SZ2Wj7/kb6Ce7r5ZEF0muuBFSv9osxYcrMRVxzDhP33QWnI4EUSw
WIcfmCL21ixOf1tr+d5LgRchsHW9aZZ+8QYn/hVg+hZQtkEzSqB71MdqTf034MIC/NZ7dU2q4zOf
8a5SpMoEE492/hi3LaK5UpRllav++1GBx1DLjyVEvqmiyjRjxV3HMOowAzPherfuv91iepX6HV/4
FbfT1hBiIT0BgjsWFY1FlGg3PlvxZrLav/ORYPBn92ZkPVX7kktfYjlFKfNwI0Zwd8jesTsWh1lg
RDsHJK4aon+WCJsFYzH5qyPbY5q+1/u3vXc0VmHpANZaRsTDnTJoCpzCM7CQMYiZhD3i5TX1b83J
4VXLcMEgyHFCK0hAFpAInG3UGad+tbtB2AC0qIG+brnElrI1QK9+zoIUUJPBhaBfbv2OdfEJ22NL
U51pQOmA+Vc1MzUIhNDGxF8scdFV9yQHYzZll6UGKPusmS/T7Jmxzxklv6npNEha0bXfb2RfZxcS
Gn/MRd3GqOZIEUPHaOVQd5pap4IjSB3ycOq1HxV6jv+g0moafcdFROXEGzJDZiY0D/4pgMytE0cB
MdmcnCFWcnr4TDAPHTTBueUw6f8b6ls5+HMycdToGFZaxxZn4dbS2PI2oSYvi8MyhiQ8xjlotFs2
15euQNPo+5hf+u6COiiM8TTKCG7C1gXlLkAyIX3UaKy3x9VGZWHemarRNz3wZ+BLBW3snwIpGlBF
AloljaBmlKJFmeJqX2nIqqDJu8dWRoRV++LkZEc9U53EJKE9kgafHsgWlaD23aQ3bGFTwxUU/BUT
OhDb+3viV6URF25DB0ugO8ZGi2/PxH8j9ZtHOUGsFScbMGZK8ksO4eu6bjZXMUVsjJizDmR6yvuJ
lSmMxG0PNRXLVzm5G3cetfuTGKYYXf7ESbSYaHNUorvZ4P8CSQ60ERfky2H5mNQMyG5WJNeQzSj5
fhyagDdB2CUsAesU3ePmYD0UZr28Dt5co1OlmNJmKqmhU9+IyMU2ZdkEfpRnoN+d90uvBiVnC26G
Afc3sx9zMZuurKP5dMm8P7NsI4xNbVAfqRlTWp/5zBonU+FG1k3R3lGWXdE5qBqtvirRnYvEXD2a
v3DuI6e98BJASCo4MeGcVypyIBl/SbsdYAFNjKS68cSTuUqp68SroyCUaEn3n+mmMssLwlPJ39zW
px0wwDn2Gu/GU5zly1lPxcqoWk+85R3BljxR/9dgvwyLPHoAXA/i+uY2wnXQ4PHA5nJGFSIRqwM3
kko8ybBkOtqbYsWYIVtpDmIQtQ45KuJMOsp1SChMJ4ZNsMan4ziZ9QixJHAu3jwmiR3wh7rprjnG
IyrE9ZhkrO6Qc4A2lGSCepz7yxc8bvg7xLZRIj0ONTpREiansUUXaUW8E+WgK9p43oXs46aSlFgf
8nk5N+ZJrA4bmr5tAMvIHyFi
`protect end_protected
