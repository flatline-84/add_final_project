-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
o7BHR3Fu31J4yZ17vcflCjVVz9nNIzyDIj9m8d1WHRh86kNn2C4sN78mnvIWmSLnycGSSccwEcLF
rECaoq5vYQ6uD+hmuFr5SlGAo8t/GLPjVsmgyjrZv6557+GRwTMwvu1APzesT/QakSusbb3l2EGn
gw5HpczuvovEyLE+VfRs2QH6MksotZRJC8o2KOroOCFRfP9kYq8OzU3ec9AwbAri4B0PnkuGZSq+
WZ4SSUnK2S4wL+un3gX66n+2GS1xMCeJdcChtd3uIs2WJXLO9iFg4B5uTcVVTsbKBq1mMOcNkXeJ
V1hCWq263kPbzopTHigOC+6PomUPMORkNigbwg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114288)
`protect data_block
DwRCNnthJlh8DEWzK8zxCgO8Cqh4ZiuHRdoAgIjVoeRhVlrU/5VbOeoYUzWrepnN2KnGp7MK+IL6
3pfWZ8m0KbdZo8r1XMVoZAXh3MriH49rLsbQIDGlDLCSTWRek6eisCHmH1b48B8xk/tDNjlbcALD
onWgMj0Jr4vBmixbniZ1ZFBHYJMn//qljICeYyfYHKGpuVhPjAwpy5SsM8ZIa7A4Q0cDfd5365uF
Xlb9RaakL26Vea1c/nDQ1JD+80DSr+M798CBn/VKk2C0X7278MWx8etk5WQyt2JBPpHlieyn0Wni
utuDTA+YhherBsARjWMQDDcEmUZIAvYgTsDNgauzJGd92/h0aYsEZes3OUzU8cjWXgbLPctN+50s
oJ/0Bj394cfiQQmsefs8a5w9dQMbe8ZS8A70GkYAQiI4JVhE6tibGZBvrfcpHXbbjoytWjqlz8ZJ
vUkAhSwPlFW4/KcVa7qsRy6iRdNmi4GuNDrr+GLrKEmzUeK7k1Tj8gxmu4W9IqFEyyE+WWMsjLpG
OiapZRaJDioGfPIpk+sTAVrGorUG6mu7fERDlDlZMX+/UwKHtTWe8rFQEUszuHIfdFAfAVTHdt5O
7XzWZMwOPt7LaFNpiTASaj1EfPQmpJG3Ly7LbnpMa1G4xuj2mUi3WUN2iLrnqRv+7C+xn823gAkh
j5QpxNFykpS2j+roY/bj1Rb2W0GAahIv67dyhyUdzw1fCzwkADGVwa774smlRix/zXGIYMVIyAEl
QsF92Cfcgi+n3b6ImhI5Oml2hk9zQbJ42/x/XrRdJlI8+fgsPwjQSfdXb+npoTna/G1CAa8v8tL0
Sbw/LKVAO7LJlAeAfhqi3VnqLL/m+AhYUYj0tdkIt4XAWaBE3+9oHC8FNbY8NW5U0TL16jf6wgSV
sSdLo28lvdojtECTtbPJXuh1Zsxarfm2nvwpVf5X/g/eKBznjlAWSEX1+EtKgfOhJVF9Mrq3Jwmy
utMr2JseRoglx0utP4MTaU7HQfvGTMdXbhg0VimmJDmngbNwTVXQHDEnRXuTSsoMQ5+OEbP08Lrq
VpNBibWir7mqon/wY2gVKaqNXMUHx88Nu1SZhtEOEk987ogrzyFd1vXRfxeA3hmH1u+37HVQIJLe
x50GeXTYLW1xJH1mRbv4ZZZhyHb+TAuV6UQHZVyvvF0s4IECyJKL4FLP7S4ylQuRIf/6gSkVY4u3
NbuKsYcSru/88qafMJcwaMt9wDARfsTVWpqhuSFGV62ZYXHuFvhN7JL3DAQ15uU8MuQ0M1mJELBr
s6sRGlDAxkqLtjpsFbR12XBIU23/SdneuJqpiuE5aZqQHarLHakYKehxSNvXGHuU3GHSegzAvlNn
1EkRg3Wsr9QY6QXLDYfDGA6vxIXLZTsMukmoayq0ji427boUqvc3fj8x+hcsI/kF7cOGMkkovoxU
xzNcyJyTmf7iJdQvvoGaVnaGgqvOLyHPrdpSvT3oJPHVlwSc+60jf5WhidHU+SFtlLDvmklvXQ8C
CF3xYvbfM5ILu8jD6RsP+EI6Awpx8p0HNZRO622N+WAyn2mKA8phnsViwGWKUrzd3+lwbvXS8kqk
r6LzJa9fHQ6JR35qgrc/DIhV0oF14KSTAIXiOoNJ7rAmJfxLohoUgmJEP2Q2t/Kp5LVBpTFD6l6S
J/fYWJjNIW3G0G1xy60IhysBRozh/nRiWMXvS3QKrQFYK6H/SdfjC9Yu1qWVj+sL/K1ZqZUf8fKQ
/tChDJfKVchK2JsJ//dL20a05B0oh+iEMMj9vdLqLFohSV5/OqXv+zONGO4PAn41W7IYkNHErMbY
h7tkt3XWblcTd0yVDBpOFJoQKtdoGCuLvx+mIDIGKHc3Y0HEcYZZDho8SZkGzUhnlp5jNV1Jrh1O
YMwK9AcXCR9o5gtW3fmanWP+HPe9dOrWxoKd670ebmRXuNh28M8PKhUJM0E68stHf9aYBfqKnniz
ds7oPI4qRNEnlWFOrO0Cp9G3FH5fJgnPBNRSNpO8D5CxiqGShhMrpJ+aujNxH07benROxkfPRbhC
nAXuDPR/yjp3+i6YCYzP3Dh6QPQXN7ysiBaYZJNR7KSMKmTEaARcIdCTUCLKG4r5bJ00NhIi72rG
ai+jgBeJ2XkPiYHU/oY7v8913y0w6VebGNySFq5vF0MP4I/btEnZS/XeKb8aXKwEFXiaII/Tlk5T
q+2WwW7tX5rf7bvmgO3mO4B1f+FRQ/36JrwHWmYvMU7AIrJGe/FFnumxQY389LrO+p/yDVP90Ddn
cEhe4Oc3FoLLUpMgzVh6o5fxyYKIN8CeY4JHsze0tOrx5jZc2mDCgsT4A/RkZILJFbp3QLIZxGmU
2hR7eBX4Rr0ObyUqiwLQWkudS52pW3ADVaJrAFan1B1AS+oS++KTDgYkcE2f0bExBn4MsXEu9+eH
64wJC0iPfiJbx60q95UiEVfyIb1+b/0eNwe+a/bqzQ5yv/CKem4AbGM59I8Sm/yI4CQ1/2YQlyMe
4HWUeIfBPI/22iQemq31FH7kchFhIGEujv0pFTYFgx4DejkHu2HTi0QRk+Agseqp9RKwjB0Qp5dd
PN+ppOwD+6yHuq+yK24CJj0X2qtYawAWEa0DP3xlNqTTliKNPtVKGWu/RzSOlT3sNX+hqmsedqLz
kZ5KqkenelS/UfpE8SwH92uLASmxWRYLMaInSITwdrLPNjdJdlGywKym5xD2kkEAMv+PXXyqlooS
RQfOkYtQJEKZkxwMfF1DpNECDhHh0b3FPLTy2TWsYzSRi2hfsYO+CB4rZ8IK3gpiB51lqCovxdzr
3yTlTG8mQ0CLi+WmMHXyGTVv8SJuz6vaQjAkQkqrDuZvl3AzAsIm0cd+fHLMTkj0+WbqDAjV8RFr
7WWXyCYLUIsM/kPxEFv7LL6E8AQ78aiim8mT4nPFspnV96FIklEEXgLeVsbBRdKul15b1pzUgxp/
HrgCdLVvlT/w5es8VTnFtQzttIk618QDU3rRuZOokxeVx1HAnYspLYdiQUKd7CSK+ZygKu8koLdl
/8vMca0AITEAYcXXE3jaI0xfSSQj4svg4EA41JYro5FopNyTrkWE7UUXUfDnhsGMBTVSbp29wUtU
jRVdsQEcQqsz8Vn6nl8po/kMdTvcS/X9Z2V1GqvmWJ4u2eENKoDM+9lvRrNVfax5vy0ROo4v3uAi
JOVq70pYXofQPPV2G6Vwbu9crK1CU1cnYoKxILAFpGV1MdXqfm1GJdUlBzsqGfFg5MyNOVaJRWl2
fi/yIka65wrAx9I+Y9nAJ4mzEqFKNsrFb342XlL/+9bQNSPZ2XLRz5wOUKbVzaRaraY0kCtXGHhg
A5Lt0n0HVjt1uRnrWRIgaRRD6R8QKVVtQp8Pqtfg2dy7QcRz4lnvasfQoT6sVfm/T2lolYZl/XH7
U0puGJ9VRjb5CSfa/2A55Ka0FrEyRkwtRbKXiRqsZao+GYtSUVTHOtFo2L05nbMTKdRf1n4gmrLL
VKUgCvaSzExPNBO01LraTErRd58Jz8/ls95svFweblKNo0EeUKU2CmWy3r0JQoVTrDgFsO4u2Qzl
KX9BOOrVTEkP+LKjaviHiSLMXLllISHkzVCGcJQwGF42u7t2L04Iy912SyP05bXjX8kOdLQb0lwf
tQlDpCsCKytEw6Sde8+Kal5UiYgYDY9vC3EkH8MHMk762eDFww0mn+xhOsoCgNOBG7QLNPJqpb4P
hWm5FxNhRoN2jGj9s8JWg9G6CdBgCCFE11qRNZdgHPRYs5lEu/lzpn1NofYoBh3seWUUuiM1BuNN
MC2N6P+yxNDyPilev1EYEeh9Jb1TUxt8J3QY8/BlaXDDCqw3C5JZbs+Br9mmpeTjPUhgjdrzSTSN
PRwbXSX9NA0oqbmOaNw+4vxqPiUuX9eBt7UUhRddblMrKQ1JFx8E4sTJOwSRbVPtqvXwcQmHaTIC
lJkp1OhuRZbnVkdN+ab0R6W6FBWj5zDxnRnspOdEyeHSWHGPUla7VyPT9M30+IQZz22q/xOIf3zj
JW9uspIaVcYc/nmRYam6BEBqZ0OmFFnWupTG4+own6/cEAakS5EviebqvbY5Wvu3BjhDmVDBMIBP
WEdeAD1udEVlpQMymxT3p+qsjxIXQVAdPi/biLXQSFuLwrMv5WDygnlVDfFh4/ZwgyGfbu0OUzLr
9CExuSCIiWyeqApzwYi38r5L51fMfWyNodP7UbglHeA91gS8YFjnmUgGSVzJZ2NfxuA2jtWL24eD
a5q2Dc96ObFT4VsAAomUBR0Ll2GMU0MUq1qD/DLGJlp5ODLMtdZ3Keqj1uNUmNrOnZBsqWL0aw6H
Cv94C5QPDoGXBzmJek3G0itX9h0qRtB64WG5As3gSisy9EPXTnThCvBG8tTaceckChGcgV0unMWy
meGibCtl4bFLtgWU588clZRk4Z1zX4iu1UFm9QBZXU67w2VE+xw9aVlZzsr4bK2VKGq8Ps3V9tJg
xyxllnyfEtEV54zqQNXgQs3moeh4DNw5MqakcRojnnN8/NEVVSyMxgPa5fZAv2vzLXgCObz9NLFQ
KHrXomW+6JNKTGX0CQTVYQ1FzJ2GiKE6uwiCMwAsJAZjRD/lu7GiE7cyBtPaKUJragpLbuKmRHV0
j7KwDuG+O6sSdN6lgB+GYY/SVVfX0V63Xqr3MihrkceRBFpQnV+v9YGWVQsaqSzZ59W/zefGJCp6
LV7c6N/p7pP4hwHXCYdIYOK5JcFvgNGsx0gcfHVWHQxDheH+JIDhhQFpv80Md3X5JB8kJ4jjtsj7
loPmQtlGgHFtHaHa4bs9rtImbgHJ7++RKuQahS2OiVKptl6iI2Ne3WD7fzvHmhdUk0BPBTUJUbF1
2FNJ9gbNH/OR15sjdGXuh6DGrxgwzyXt2BD14xGznGF7QLFgSmEnCzoloAxM+ujwAP8dVFoin/GS
b8zmzs5EoUI4NfAlJ4Vnx1XGtqTCb3rlSbsPaCs1gHy41yWEyimr/bfgdPhLLcVlUklI5myZ14OW
Ep6Q2nn3Eq8Qcw0e4Lzzl/3EeIZjnrid6FWlXhMmK4Bvj+ddd63P4MoRONv3KBL7BAqMQb2NwJiR
ZodD28CI4Tnjj3WpWprTzIcbbOp6TxvG79F5bcsYgq4ZarsZMzC5IHndoAOLmOWe+62geKN/68AB
ZTjpVcU4+ebhx8kDMVKgFJhV00F/341k7DafzRkQTbUZ8C+1fNxt8IR7KX5IXGDO7HcKpbmDaMJP
/Bht24jlyQrsu5W+ImO15v4rWBt4PZiZuAHsN9WLIWI5D7INQG7GcqnUcSPuy3FSFEfr2CvATSJw
PGeW6gzSAfe5+CiHbyHQFTFZrZ2jsvnpjRPYjCsNci2vztlqd0p6YfNOjbY88luXph4Ey0qIkjbZ
iEXc4HxjvIcvETXUM4/v9no50jiE4nrbyNlZOF5+MdahXfMgYglA+R83GSE5XHFG26+ZRIqim9cs
4XjyenNVcAqzlopN3uiFKCP6miGkoLqSvuk/UQNX6mh3GSv++Ii6xiQuzqDnXTbQqLiMgioEdYeZ
M1ypMxJY6+fxH5qktUC3pZ0phSElvPwsdFL92gJY5JizC03R/v2FmxierBps8uxzo8RO8bQwqauQ
3B4ioZZejsaO8PigLe1bvlSOU+UvlsUid9+5kFsMslba9mMwFfupVLl+Eh5w51nJ0jn2vzKD3M2b
qRi5Y71g7GwMDDRR+GWRDhfUgx5dHqtZyQFUC1qVAJvXtyo3kkvUWv70shH4Gob3SslMdwiBjxwA
p1nVaCNmpszMHD9V+DjUe2lHusi/YHbMN8EN5xdBiG+xL9TQuqUIlKxWFhNHrVTGesju3CD4Zdkt
IVC2VVLT6EHB048a0zfIlUhT4cXwB+3LIrLGe2Rkab0h99io8qfv8re4lLr9Cl15hybA9QlKaSgN
G5d2hFDu/glNjIgNJk0yiv+/UuJmU3TxM7ypJeoxYKbGYrMcImoH3hjDmrCona0Xb1xC2kEDKjrG
rxR41/OiDhKv3EiDCNdNVxRoduBe2TwYTiUsXb7/IMXZFpJM2xB60skIsXKfbEwvcclDdcx33GEq
qsHoPWZmcyBxeb8wlvn85zuv4k29hnAQXLU2w5oTi3owZ5ecWFE38N9om05h+n1cyQdJ44tW/Au5
j/zZKIs9/sjrMTHMxX9YvNpvHGAM8aayUnbrdkzCNi/oPE0TBoqGS7aE+oGM7F1Lk4BBvGRumzMD
nVeB+UYz3hR3nQVYBQ361RorHcqz3L3KFGd44whANxSWnVmhi2ACJ3KzKg90UA4UZ2oLpXy//p9T
ziL0+RHoXsOWwDaTYu6UFAycfTSF9opPjB/kvi56gU2YMajmttUxXHhWBgSn2a2EscFHN4KPlXTt
40l4X73DECoWkwFTwVKpLXcSKliB7ILVlsQ+BSu8s/0wQmyWRc1kaQjXKqaQ/geigfmCtP/iDLHj
7VRLAc160Ny4lfwPnzRPHRWBrJHtbEnntIQu7ww9zCeN+MRNNm3kcdmwIxnlnKOh2MtG1rKMPhsO
1SMzGv/ubjZp34UaO53ByCVShWi+7NJd6jGYDkOyLGSf1tlobj5vBi3cm8i20RqiMmttX62QvAuR
qWvXVB/7vuV8SVC4xPT4wQradgAjHWWzTxGC+hNi4orgpZcB3v+Vr4Qq6FnuT6wXMZ3NYKTyd8dC
Wsjh6vrorYbIOl5n1gdtJV+BBn+OU9n9nlfHNO3vmarQmuxBTfegBZeTT28uh2N9k/kNzPsXGMd1
jsIU9fL2oYnZdwsdefiIoWKduAiEMGeLr+w3urK2C7k5poeR6S181PzTSDbLMmKrmvZf1wZHoVuF
BpXerJucsoMJBdTe3/Q4g1Jjhh/duk4tJEzd2uG5GGHizBx4G2dBpzOlOadUt7UQbZt+JRTJOkFm
0hlAaKQJ8V62Td9HvwuMw8gwQ1TQGfCG359hV+mGNSIV9oOFsKM7G6froae6wX5LWsTU0tD4CZN0
7L77fY1N+1L5Bjg3r48aPNU45RmXbfd0UsoqPCohiJalkRcwJ2Pw3kSQ2nRj2DFbcDHmeO2O7whJ
2mFMb4bxDvQXFRHSIyLmtnY5JL7MKBY8EmL3nfNy3i7jO/hqWLslNCAuglrXC2Vi8H1hc8Y+1Tfk
fFWLYBuJm7sQ/fWKyBNpZQaBsAsp2tNzTXc71B/hnvuM+qvW9XlBZJOAdZhPorAK59gAg0cikYam
s2Hxp3q/g3cfl9ukN6gEklYpVI+wzzffoaN5GiTNQXmsuVbVNhvKVamgjHyouiXzO1S8lAYMW21L
3oB/HQzq5DRn/Y44nzeS1EFmtlyywIxJnRjqsiP8Rh4H51TOfxc1fJpbQjMq7udjFsGWVeIHXrRH
U4KnpFVgCS4X9Gkj4F7UoBgkC9usg9Q7aT1pi1iEb5B+uRx0TK/6DzCbnWksKNUtsyiAgqW6kunB
g2juBVOSiq0ZAXbSBU2Gq9zpjYyZTEcG774ZrsCAUaN0ldymQ1bQ0yMeL0T6msYJfSv7JiK/8r8t
CMzBTqc4JqI38T9xlM0ThVM9OSuN/fYazsVO5aN/rIVRlPOIMla6npCJo48SctWv8cuz5blIdW3G
V6ANyuv5RC1mWpXbvd792bPYHBiqU4fPmd0FkV7THRF9ety6JWzZAbSyOgawYJOoWfS1iE7dDbth
pnUICeyTSpu3DPp8jJy8xLJczBiGi5T3qwMZLKL8Hx5ggCTg/1RqegEUwZBibbCgCc66JZSINGad
/FLjCshA2wHpMPEwd3c77Aa6euyzy45WtkdRXSQwmr3ju3atiTAoMmraw8ZPW3ERh0HAjTr+a9UY
9sTwQN+fg39RPlseOgMCoit6hJLn5++SQWIFYK6tQgBYRA94X8YUBQGhpEU+zKT6D+whCCGNDk05
jdQD0SgJs2FJjqfCy06FtyzRCbJqHle+/iL8ialsgq10YLd1Euk6TzI++XOnSfuGD2PKxdpvYxgV
jIzrH5J9+BWEDt95qhi2b9+uPF99C+DBq/JX8zwZg20OoFaE+vcFwOwPIS3UYT9Nheel23vhooFk
DNUFu5rmLiybcFunzAVteOB5fAEoW3df6Ei/gIhIqAJfoME9XOhkQFLdmEmxbKNKrcMLCTman5mm
dcbwrlDUEvTHD42VvvNw8E7WQp1QEv3LWNxT9NAt5z6ATYXj+/3kUJFRuFQpSVAlw5zcs+0lQDQ1
NUSq6Ll7fKgDrzjPsKdQoDZhZr825ZLCBA+KN/84fceMV7LbGikAy4n9nBG6WlVVqBXdnwIgwFA2
cAwzF/7qNAk08wVrIE9OVji8EDplm9TInejdf97X8P0VE2MnzfZloexDbgZxn0F/ozNVcpNp7edy
OvMaZfN6Pg8SUuJHoMg9tPc8LhuvjL7UoPnVebKAa+Bs9IljBS46F1ycupjLCyAql4d3sg8RdtLp
DSVaiTUejPsgfrbJKi/pXMtsQIIf6FSgvnnFsKvw9/8iW8+GA3L76B8z9nXLdo6gVq1UDFeCnmz5
RO576/3HD2H7hU5qpVpFr2IDvdZeDHLHLHnG1ys6bMhxgvpwonfo2lPqjEJw3FGwfUVBbgqk9Ehc
3ZZ8A5PA3Gb6QybJy5G7OoJQ95vBd0OfVs5TSTvzPZVWWKOe2S/+ad56pcZOjOo3JI8IuIElEGw6
WMzfl/mVunnktNSFYlbwSR60JsqFcmgfau1WG8SIwstpqSIx67ODjro5pwPgBW2po1pwMAyPi7Pr
Rb4pybCcVzOfUbDi7TJysg1NOqYt6pW7mIHkHhwr1fnpvIM6q4EFYaId9jzoAOgsjJgoWvqtJxkm
GqJuFErDTr1/0IqEVn9iCtrv3YJrAos2V3y6S3G7iP4KbXM0tzWxmJvIFIP0SSw85c6EkkZWdtaF
HiqxhmteKiSCQQ9bs7MDdzdTtnc5xuJ4YcOk42Z2fm6aFUMlG/EkPmEBbDLN5lm7vIkQR9Q5P6x1
IH/LGj/ZlHo2TUN1ZVirRkAFRJWkfSPkiDkbDTklhxM9lgKdBqWdQ5m+Kz4bQjUhNyzTrP2MesmZ
erx55566IlA80IAmFynWFJUvT37G74jWDKa98GJG49P74tgKb6HS6FXvUbLwvhV0RP8N8WfLRJdJ
XWJg/3xK2PRKTE5nSAqJQgFfIeWSJCP+9CP2IL+h82v9zGqgcRN4cTo2jF5rPAruzoWxfy12aNc2
+HnL2E8gMAHvfL/qzT7zbltlhAbyrKLyR8vKrXcwB3+I+IfswF3Ol4ewLQdxkzbu7+eqdWk3RnBB
/TKFXvCy7o68TyTeQpIvf407e06cVFm/oz+yGYiD0Xm0etx77+IyFHJVh7lg1Wi369rDhhKdku0v
tZFgg89Hq4egsgnLko1KuCZ2a+3Yji7k9vRYr5w2C8V9n7gi32ht5AZLZ9GdS6dwCpimCHtXKocw
TH9sbuTSFyN2vjL4IUYcb29YaJ3dMc6wIytboHfT0wNSH1CswIVU2QB4y9k1dj/ulAl7IMDXSyGn
aENNuLMtc8VqvaE8LEJ5+9hZQCywCJcpLstqubUNFDBmZ9WuCrG9bFKKBlTLyKeP9KAM2akPlQ4J
vzliSwZlRf1m6AsGJGtQm0kXU5umYSFVuQn35YcaeQNvRiiEm7JDSBvonPMU8TpuHn7rpK8KHURv
2f7XF20EqiNwx8QsV7nJb6+C5UJ0W2zCxI5TX5apJjn2eGGrk0jruqI014mNGhB9ZgrKOALyr7ID
MsiPP4YEiWK/wHv6HfZIKUA0AVrM1SOwa5tOOA/dKNyrGoZd5d6C+co5fHpKQp2XDSFh6YbqUtyd
qY6ZeIUyy+F2uLLFVLUZGZVgMIFVe5xme1IdisgMVQlCxvv8eKrKnZguMWNJusFGsmZXzQ1UHnb4
kcAM0swzI3eZNoe3mbMS0hNFnS9roMkBDTuiPfByoiv3XGWVl0y8LBVKZySTIyrRbdmzL73RtRVE
lI6dJMKusoFiHXi4/b8K4j5JttmuSV27xEkariL2iDOjC2KXLj61KgBls3gd/6sz9HPSzvVGq5Hf
0H07QZUkOkVOEsyRu7BwUk0VfKnEOjckWlp6wxxMBCeoRoxOjVOpmkJdc71dsNbwZWmK6qBYos1W
lH0aKQJNtqvw8x2imj/ujhdz9B27+9W+qdz+3q7r1XWTKF8ayFfzmlFld2aR+RQv+4updIzCYSd/
uWG6/CSCHpA4YxqM0RjNxVkz+lG3XnQXgGLOelILsY1eI2A0fpOfTEHL7igpnZqFkc088S0VMr7g
jKlxBRbVZIM8LsZJWuKcpakXEEwbnKXLF63ApUVz0+nKDX3B8D3ivty3j7WjSaLHfrNkbTYUeItR
AFwhoI/RYp18o7b0wRbGXTwGiJIFBiMHKy67Xc9l8L/yEWy/EZ8pPJqPzoZqk2scWF57NXm9PXjF
CyVJGe26S6nN3aRYTgXVZojBUd7umvEDaFBQ6vqU8ySJnZc2GikkFoqYupDkQpnQKfAnoSnLt6nr
03qL/pg5pxXVNIxvaLa5CAvWWxU++lOAT7Zj32T/wsRGTUDjgtJJCWnn5a1X3UvgUZ9+9qUVe5Sd
1DYLYrkw7/eoECpXezU46BERCd6Rg25n32Xu4/CPEc8hcKj3oFLX0QBKE1kZ3Mo5lQVByG+JnNYF
zNJkPT/vDCiq4o45N7BjaG2GE2loVO6JlOGhp+KWkBCZxSwroDQ9qkluSMK9j6/TGpR6Z7brZ1uC
doRGu0jVFy7sy/gXkgK2kvdP2xoPaA/CGwH3a5ew2Mp50oTnpfKuhSGCevB1Lgc8Uji3nO9cgrnG
xpl+gNSRubz8mxqIjswLpag+cisAn+Zc96CYQYK608GsKlOyoituUPU1lTQiW7Yyh/bINDQrKW2U
1O1WnATptWazLcpTtw9D2IuS+k2kdv93nTB/ka1FiEXs5FPpycljrXJRdNfcBflxqa7vf57F4gpb
ro+WXJj0JOWyvNjCwzQoPXfTqRJWCFOSZy6DEPLJ9OKLrB01/3lw2a6wWzRy/XCltYPbPX8BVNSf
eOuze7eLkmjNE1VEPEqbr6BH7zDjY86827UVGDTN7vwdP4G/6TP+UqslAvTuMnJM43ZQAf4eVWr5
g7GInwAd8Jfe0eiXYkzzcMSkWH2gifwY/S7SVFDDB7zAcUl+IiO315osRBg5MjB7bDVxtBhu36Gb
pugAUprwAab/9tVhC1Dbcb4Ajv1gDNou1dWWmkFjXuZj+raUtHh7DmdmnD7N6vbLlEe3+yQ5VXvg
mROmx2p4eVJ2/fNMXLIGcQaEinULEkbfyvi9jswQ4D4jVe8xL10mvzWyt+0xVCXt07Zhshxo58B5
vPrVc9X7Po38XOqIZY58M17Auy7nUZEKOs2QGJn+vRQOQrhlItDyAOefKyfkYh3GBuN+Nk4VMuUy
7Jn2EyDNgedshmkAj1qU78HAmdlOrlmWCOWyYB0gXlZEPj25ffiMeTyHK2DsAeT3jsjTUJLbVjcN
aBWhYxT35+tMA4Nb0n7xUItjTCFjJorPLCbCpoDlhgr2s1fdAlGm8XoswH1mBpL0y8ughWXkYDes
YpwsWQhxqYhK3Lip4xqqZ4+5Vj/dek43GKz3/qRH9rph/k1LGRbkqbbFmcwm3qMdRZhKtp+LwR1/
/Bdn0980H+D3rnKJ9zN7LEgil38VPnv5mGxU2Ay2bfeOiw3T7VV/QnIVEk2tUEpFZxvR1VSS7Wgr
iLlJrX7l8tbB8xbbXwe041fXvH9btZwjNuR2uhqaTFgAHXdGaH61Pj750p8PNLN0PmT6D1TFb5R9
LmBUm+iFfRYxFaOVLPv5jj0mVaFfYrwfINRpWaSWXxbebeUH5/BJpJ3U8TD6SfTr1V/+DERj5Id4
G2UjyclPGEVnPC7ZqqjZlZL5Dq85XcDj695yjn8U035M9VFBPkjiXFAXmDyIBf0EtXmFzTVgXvbJ
23twAqtkJvG6UqBJMjx4ZSfmC3zhgVLHhRsCJU753dhg1iiiEn4dyvzNFLaxN5XjJtqBnYbBtXgt
UL+fXKQG64qzGJjAJ0iOdJSMKTqdnWTbf1m2g9i8CNMjdAJH2zFCSAOQcjA/BwxAERjb60mUDqgd
ACJurEGh/xu/TvR3YKwUivUYjzGjesdDTFLaPcol1S+B6uhAJFGndJDrgtL8I/enyPH/G7fccEAn
KJ0m6fjBoeigoVBU98xyQuI1R7hBb7c9uVjLnVbZ391WvzpemuONV4Xna6DUud5tHhkqwItT+Pb1
gDde2/oLzQ7bpB2p6RzNSo0UBaLCvDGatKlqynO5lc6syITLfCIPbJzJ1by3vjqUF7olEC/engOb
BtDSYG+e+gTuch7iL5mUhK4g4/sRkPicRe1piI8Q8BikKhMrkTG+C2ndOnZwR405bGNxIf3YUdB1
9N3kC77URpdkfpBO6amS2QyX5cn2fIPte6fHs+JIRIlU2F35jj3tSeig4/PPu7U+lQthE12L+reA
WQ5zMMrlKsg8AWRiCN5GgbBH5Y7jf7M6VcTadT8pThe3EzDLZ/IvzhmBuQuFNHcNsehsCqmwMXN9
1+QUooY+xHH1Qt7zIOekdO8AIOh6VIjlA38DHRRVs6bJUU1ccHqeW0f3rskF8ozxqx1SwOd7h4QY
P4bTZKi5k+AYNCVLFm04MS3YzT+d/6uRc2ywFzSXUPCqdFWEGeF11w3opyxllVQVrbtvRNtu5t4Y
jvHxRFEuvsiLypqoJ3frXEaom5CGKbeJkeftHG3Iu1p6p9oslrrmL3KCiqlCv+5vS68YApb0TI0u
enoxxdrY4/sEe4EoIwsG8aWGujATGp07dwVBd9loWQZnMhjSY5OUVu5DPJhT8wlFdMDcXyvaX/Qf
A0gv3/ovRP0VmFsWforoJtPJLgQCXN52aDNpfUBjNam8j/IZU36tEzVNt+3FjK5K5LS1pQ1CO3YM
ZuttCTUNqj4hnaUa475TAJ1UVWUc8Eb+k+I63dwITEebrtQzWrocE3/4wUo9edzQbTzWsvR8Psz9
2dSL4lDqh0+8ZblpvsZveB2gYLwb4ZRovuxcTho3NXFm+eyEOxXua9/NyRfWYut0OhdM7k999BWE
3x5eK+bfNdFeUfIY3bHg8ChLyuAxJr0vSep5SK4sHI868oTNX3maozMXABtiu0nD7Qt6AIICdJo3
pGILFKehJP7+b+3NjnKRe8oqbx8HoftwgXiV6y8AanRHbWqePHFeYxWTlbRc6y7CBBxj4o6UcdZE
BHpiHuagegFpX6nV0bBTEDG7Fu0GqXften21x/tV0ACkMQ2Z9Ycuwp3b2GSyuSyBXQAw9SmI7IXk
FWRNrQoCIpMqF40FWOj+iEMVEUx0GJ51srmlGJG13ufhJMBc1DyxhwF89BI/YVF6AmyKS3wlaU0T
A5GCEWTaZamZyDqxmDfjcrgVr2tO4YR8styZzElewMPUwCwnOrflDorobhgRo1jQREWV8CBFKlLb
tiezb1lkLGozHCRKnEOmAeoC78h7htXVXDx4pziBNMNTwHwGQ1+iub5v5MWtojwQjJ9zE3M++Kxj
eF0zfPQJz29vUeB+4g5v0VBXBB9zTqxBGPV+jmFRmKxfook1KQaKyfEgOYNMeOqtRL5zbR4EHVse
eedceMSgoxDG5+c9CtaKWEO8+mm+fcMDZA2YHnkb6AtjXe3rZhx+MvRi5gjrFo7LD1ik+63gxb2y
A5kiQHdoPhj1PkI/8hDe7t6yWR9tVedPmNYL1GP0LnkbCR03tDqLPMCKUzz7zFIxidJHtvf7UNd+
P87naOuoNIAs9CX+31wAekeyb8KDSjtHGUAqeZgiqyJBDhl4Fz6l7uo4sXjrtVlHS1jujCNnNT/p
ba2DQTtBxZJzw6fdJCKXl/45xT0XrZT48n7TISt6cmJIfMNu7i2pBO0BtdLiav4wqzOWOQGChH0A
tRQnj+Hnu0ugRHITOXMjJ4v+d92g2nL034nrMAbGQeljpuYgjzt94kANaFqmW3j0TkPX4HlEvfx+
kKose3Gm1nk74fjmArk09KKpiXIUIti2sbb3Kg6g0XJbO61vrYOjR3bSSwZjjZ6I3deVX6bFxa/a
EKufnzQVtlRlAcsG7XqSzVhDREAsk9h6rzgY42Nd84HDFtqEgI1RVTSjimnJt2Sxi78+L/NiDwuA
lv6oteflpqXdNjGX4yN2eJuBzwVbkhRbTHwbhYGg5Md3fZdc5dhBUHvetMFq0jtz1YokWxpHR9nh
MGNTz5l5K2h3ZiAXg52ktDDBpCuJkCIVu+E6pymOrUyS8QFQFb8tNraWUr9nqn3n/Vg8tjkorX2+
BYJGpMC4CB+zCPmqTdef3VFfbLQg8Sfw7JmNqnybkiN7eBEv3zv7JFVZbJVxg3kxqwhZykguCi+K
4AiUtGCAwCjvZNYzKKCsiAeO+wEPfx0SbJeVih3OcfP7b1lCWGVLjJC5jLAx5y7yNjnndfGCke1S
TZx3jifiVGBmKxadSXtfSr4hPi7P6dWq/BRHSvBumzSlVopNSymBMV0ujw6IQndtLGAVJjoy821i
DGrNW4uad1SG9ulFL/2eg6HvbHlOMXbhpjPeFSyqrsPfvXxMoQjxuxF4yZfOqJSVKPK9wvs0corj
Bythu92P2pieOTR5FNUzLAZPU37bb9ZAOEEKYZ93Ilp/j5JaV9bqZoUbqxDIpwW7a6GDAAWfphXg
Kf9uxuGN15hUfwGal/xbE7sc6etRX5ogjF+jHgEQBcrG32OIX+gSRUue1suGSH8vkPphMe+DkNy8
U+4YYnGEXH/JIKExjNhMt/4jmhAvNF0tQHMjN4WW8CW0828kK/P/crqosiGAiRfmcp5I/KojiAUd
XONV/Z0HsV4Mip80KoygiJ9VlWMwXem7whg4iHBal7ugqdJZ4rDSR9JT0wu/5oKcAFpn5hZ95W/N
T8+plJzdVfaYulelGg1db/3/pXkHxq8CindweMylR9qF2+fP/YYkQk77RkhlYKpjjPdl2Nshb+yp
6/+2qq+ZKpXYFAfawNSqIfMEzealnw8vDoxizfryqc+RxApz12N8D0qosxVvAX9/ra5x/NztbpwM
QFkVY3iOMBNPadm4MgunEOcLhzfc+CaJpihOiB99lOJMoyBA+VFprSGDwsS+L9C8WMDwfTu+9KnV
278Y3mncKvXevtK/I+d59cVsmTT5/TEluiSIH7jdV1I3PY9ZedNu09ybWJYCTh0uz53nWFqBHNHZ
v+Bl58dgDjOR+XvdkFDOFZwxQFv133toGA+5TrNvnXMtDaORe7Wvko2zNpNh5r9NTOkvcTqXr9hR
6n9K5VFUuDqeyP5PgZEVHcMz6dyaf6kAhY1SawuhaKbbvaj9Xjvt2GUv7yB67/oU/hnC2E2rttiL
/90l5V90wCGGn59AqbJFAAkO71ipmRXFr2dDA7Bryony6GcgedhPRnyBizqI1KGkB1ciDzHyy2F4
HhEkH8PXkFKB2pnZAVClhAstUtfSq1IqXFoWYJu0feUsHh3sAdFPHY5RHGN5SGPL+JoRFGG0V4c5
ysRek3NHSiluncqe8Omo5829+gRoPsyWQxjMtU49kuTK2NGF1volQKURSbqyrd2U1hABrRYYQAne
oLVNPSuCVswonk72sW+fpAaRfPTHWoSizs/BiAVKs8BywvIJhl0CBBD0rTmcaRnnhqWowSwPV5lB
kNoKprmHieEqVBpEufV5bNq11YMnyddVT9pBbVveFGq+S/17ExyGAi7Iwq6N2jWW9m7VP5iV3ULL
mh41wcNHpszVhsM28XgRlF5t60zjPxuV5GbENLeew9AMRcUkrt9Smu9CtoIjhKgtv02f4d2MULuM
sbb9PZiwuE7Z15nNEfuu6C4E+DscwD2w8CTfWb4lS9ozlMhRIDoXktMRgZTOSpXhn+KSGmV8lYvh
f8V9TOl1TJZscEoe96SP/FdZZphvLXuotYKFwgJRL24D328rHNl8ZKgP+TO+5G1t0TIZoD+uG5PT
se7kEehaYfuMxlsQcom/CmziSMrlOSjEtjnVA1CHopVYTXxyF+1+LPR5aoqvAo66CmMdmLogNrm1
as/pakcfd/eTnYtsHSsCv6P9e2t9tb4Rxs1Z4salYWsTL+7VFluSmLZXxhMwxMNnjF27PKSyziSj
KU1d2GKQ2mOH4iw2EDOkJhPggOJdUv0KF0+g0IFrB0F1FHf68CPCy+gOzibE9uu4P4blYJHgjCWu
DAfYMl0ghlrkTMDrSK0n0kapooM+BfW3X58amoLz/wZUc/LvVvmioYA+2Z88gtKOY0iN9ZFzNmD4
p0pHJ3WrM525zerOUGg+fGKHO/RwLOzQrwb5wQg2PopagmRWe/oCAfXaKBv+VOEjBROTJXLDnBz2
mbsk6BYZl7VC+x1ohlZ6zTtuWnJPd+UlAP7zO//aW9WDviShhie4C9v6C8Zh2jEsBM0vnpeJYBxx
8urc2533XsQCuw6SqB6QiQYJniGjMgQUahmJhKw+BU3LJiE3lRIpDZ5b5zKWuxmrO7MidYfFnz6O
O0P/HDQViDbEuzXb//1n2KdLs9Kx+4N9BZHAlSbaxEeZDiJGwXHGkxGuC4Bl2ww8h0br1wcYAels
GRIg2rfnk0csjS99+3a+guTIunUjm28CfBxqSxC07dRs4+YSWkjA+9t03d7R8S+zZAdkRr/XF0E4
yOZJhmXtw58vupoFUU5ys+ypDKbXa+lj4m2MP+ub+YleX8gDAHjp2spe3Xpd+oaCE4/xZX58yDCo
dGZgUrxtLqc9KTMmNWeR/9SZBAj71u9wP4xQ81AaI56mOL4yZjEqFagXW65MJdTnk4aPLmtbVI+7
+g7zBjwQOUcCORdFRD8xQZdICERGSe4eNKTHj0O5efnNREJLHDxtCFOOFLT8U+a/P7ko5R8/SrJO
Oo4DGTK7OedBQQSbocXUmSIixUZqke8tJQLUsJDouplrpWJG0u1XFJJMuhPQTgOC+iQLysonW2BF
dbrQc5E8gCugNcrCtV6h4tgoBH4Ai+XQ3FXELe69fVvSN0ZGKksl1bUE8L2fEKOqYox0M50lIcze
bt1JsL9Ku5XnrMS0RCevZNWIkvRZ+OwWNmkRnSKTQknjhgfvPk73Qhd9XH6yVHlF9SEofSj17P9n
vsACkr0vpTO2sH/RL3HLw6CJ+rDuSiJzYSWBMaFQjtwGAkcP6UM63q5eIo4CCCFNwTL2ISwLHmsx
uintt+I06Lm7QJyveg/+NKu3DqGWqfN1C9aWMzcjDt/8rs/gDLkO81SRty87NqLlIlIgoi7pcgMi
jqsKD8Nk3rVBdVOvqX2rFmOYfDCsNOHWFUeDx8q32OgyFkSUVGI0TY1QgAtcGItX0tQCQnaoTt6g
q22h9Mc+TRmp+pJEhXd+32vecfqEUDElq3AoTL4VaOn7il7t9VOZKvdx1ZTT5p2yYIMGHYARWOKv
hctn+PYFndSL+AfjCKyUdAWt64Q8CJemc2vi71llTdQoVlCrlO7VxLTR5geknbGGRTM51MMeGNYV
qcmGx4fu+x9sTeqgfcufUtPiNuHfgaH082IDtcBPaJmZ59MXvdMHrqs7cPanzYCQtaU6XoxVDP6a
uBUOXpuD6uZ+C87AtyCagX3mBsngqKr1CNB4Bmz+UOcxuoOClPY+SIN9Zk5wHiyM8cHY5/0MptfM
E2B/ZVVJJsZjPswXI9PyDuzyeImgz7T3oWlVqBM1qkalxTK6cbCJGbb4ZRV9cGv8++VqGXwfE6CI
9iYPPYKJXJKfVEXIah+eu9pto1rKxFQWUHXC326U9/dT8bj9tdIstradD6bHggBcFxi+5VwqEj1Z
aaNHIXaLr34+2tNToqNFTnW9P17U5o2YaTNP96Sjk6vO1JgnSiobhmx1CcEADeT73lhR71gzJy7z
HqmY4bunUref/gK0rH/HlufXeYn4H0/CWX245SnaRrxSNYC3wd8CxWqYB50nXD1rHijpzEzvYTJK
vQkTGGNOYyNofS0inLdlbeV/tV/ESsZeA8wDUIMWzQYo1/ZNndIQ6a7DAEonS7zs0redbVcc2hH7
T5H+T7nQ1vWDlYnPDihasRlNB2bK67nT78PIWYw+Hdcb/K+yJ9gvpR24IG/9rMp8bUTNz16WvAT8
vl+oEff1Hq597Yd7vmtxg+8zWloNx6CGM57uEue27i9J/MpeaZBinkO8hgOf9PRpRR4/GuXeYTGU
LL1Pna5jaBZSX6gI9xcHJMB81g46np4XP08sgbA4iKHcUOVfUJ13CJAzzi7UcaekwmRjP8NuQXIo
csTPX0je1/ajjyf3i04YxCzy2LFkBdQdGpDJVM29WvZLSvfbePijZ2gcRZSxjuJj/uSFr4ZZ/1bH
6Gq/bBcnp18HMtn4UafxzwYWYlOXKJyItOv1DSL8hu0c+SVaRqJ7p/HKQ5SGeBgxpFomqaESOkS7
OIaK8eSyx+aqbdH//TQIeS/ImvKNaeNXf+emWnLJaZH0zBFiBjUOMS/YWS4aPa/nhJq1D0kwY5ZK
+eBTN8ldhWcB7Q0wPV4l+aGa9ndoBPqmRnqy2KW0lcfAik2Dd2db5StGms3/pJSS3VO0wcyp3/bm
fwQBEIb/yQRI0flXI23Q4ul+IletvLPLjV6qrJ8gJsOayhuHo861EQopQvcs4XvpuKBVqiw21dUf
WbhXegBZ0mGlSL3NKTcNdBju3o/mLuOoO4/0HzaRzEpzjX5tljOSDrm2Yt2wun57JHNv6KlNr0Zj
TAQAPRTGrMzNJUDwDktVUcHUnAit6UN/QYHmpQ8SkWF+EY4W1MieEgg6WDy8bK0Fv/MIPJJTew6g
SFh7TY+wfHHSORaprTG2tZ0EC7J1rWnob2vGP6YMDAgeQo88jSqMEbXiBmum9h/kVwAWXbLkdRlc
3M4LGFj+0jKSmFNiXIkzW85/whjJCMMMToM2KKTRuy51WkCZe/RTfwghwk4iRoEh2Hg6i7jR8A/b
9T2ld5hZ908Rljm5yc9bXS45HWJZAtr6bjDVXRG73lO4Qx3M/smEpuYpoXS0vTkUr1F/ll4bMuRu
pcYS2shKCmrS6vwuKyPEWMzTG2NXA2K+wCtpiahBw9HHXwu4b0edEQznNGopuN+gADAl9cCPI9Uw
D321V8t0L7YOPUeRAW+cGWO6c4fcZBwu5DtQtt8qvkz9iRkPcLXQLyMUPJV4ECF1eqhIia0lz4Mx
FGXcm17fnV6ozD8tx2z7gf7ZzplZLMdEyhFUYbUzW7KTAxEX2HKL//x3+GbWMDqxxHD0EZ05QmAh
0iYIsfI85nTG4ajF9kxgmjbkEVwUJEb7jte4KaiA5hFaOv7NtfypnkP6otg7sxHCgB6yPY7kcRW5
6JPtBw8fsebMNwqY1nBXSEfb17uqxszHG+tesJdhPSZGsMQteIxYVSOILniPDKy+vVGfkUM7enGy
6O8Q93WIvtgUMgCD0juNUjtRG1sOwgrFFnciborceMDqDop5EJQmpHliLRdyMpV6VlkJrBiUlV6n
FZlHcitcT+2pSdmhmbu7Ks/TAZbATvPTTga17F2Xo/bPjVXAfcLwqpDWR2mSRfhCJ36t521M1xvm
XFaaNl+n6wWsVQV17+QmzBGwAFQjbzig6NS2kHCgLhG/hEpjtO7z/gUZqtg7U2UOKITmHqlKV1PF
EI+YnNYya04EP7MzT4QYYoFqXIdSFUokBazDKwCkLl3Sch52WKPR2n5+ampUeuXPeFrDFNy3m3QX
dHFQo9wjsp1Mv8rQvYDpOg3Yrq/IBgpZx6P3tAYcgRDJQLo2K1Co2sqUGqQsd7SCf6oG5FDnRn4L
QYBOHCHpRjD+03Q/uWA9+/ZU89Pus4cFeXCJngvJ0/mHbpCMkXemol8eUeuT9O2/XYhf9mauJxPn
IggUEdVdk1hwTxvL4dbBqAZlUyTRvO3TqdMIQA87j+h9/rrgActAA4yF2Pfk069PnCUNs2jEO2Qr
B4zogJEReH+FkSYbd6gVWIOAkzV+6RdlN9sCSkLd8rHV+W8yx5DeVEWx+0C6bTGiPvd5RbTGKm/h
t8pVfUHAPdn58E+Lbn2BsvlGI0YoSotdNa0AclqkEFuS8VUEDreirKy3NUMGZfBrZFI4SogfByWn
vq5B43+6T0lb14X5nYyvb3PRN3LL7udrK4OeUJU/mqYhVTEtV6s494P8mbl9wCxt3USAvfdBsxqO
EfJfqc+ACKC2O2JGJjaYLU6JIN6vqWjaXw/YDKsrWqCONxeWOtj5AoJxB1Rd2QUp80jAbOpdnjRw
IhgeMG2/gVy4b5tgyES87CTBjQxAlPKNENYfSBsczFmkAhdXH6Xw2pqpQew8IV5nFQ89kbQoL2rX
MEVRM1mhAfpsxcp7JbhMKaglXeqvMKjyxEQkaA8kINIu/M+lG7uhxLgvDrkmtSpu+tT+cSGh+SrX
K3Hhso+MBbf/dqQarPNwymjcOmIRfJe0nKJtpxS0GFU7iw0c+Q57829iVgSukVkbSPU8BHN6LDYe
DdmHjjQTlyYN7mYKWyINvWP4mX1di9huJnSvLZsilJ8A6BmLl7ucluVOZ3duZLL2Iprd1kPnJEIN
LnSI7idXCKeBhYtDgaV/VgzB0reE197RGmLjOaWj8C+QB+PwG/BnydRYvdOAmPzL0qfY+Ym7SMRU
Wh6O+jDBwHmbTt5qsJNaB8t8YhWhO6tBPsEF2iUihdtf3+tv8T8Oe1ncjGwZRV3M/ddwDxdod+bO
ZRsAX153kOMACSYVSbB/BOXcpyZIy/o+rvW4AG6dnO6cnP/LZpbxPycXqqNgd6c9aDnqQQqV+nWl
Dq+gRPZJjLwehdshnDPnfDWKW3MS+vFFTbbKO2c5FuWfHVpdQNqb8yoyjxqjCTYOloeD0pjijpLi
0pUDSykYABWw3Ayri2yGrQB9JXTJuEYBH4WLtaDczZTJzhBf0CQ4DibvX0w2ls0B872yypU86tP6
XcOvsszioTqWQfsf/6aMN//YiWyIbt/ggOyyoT/f1aW4c7tXB1r3bvxRvJ4OibDImvt8c8vvU3rc
uNmMzRV1V8AyxOfsqCG/S65PRW+SYk4p0pwLG9k063dl69235AnhE1qpo5ospOh511+GBJnbKtU+
5o5+7YdEmvdTj9CLShOSM7u5/8ErZZFRtna02XEIAmKI0pOfGQ254UH7ohekOpAam1eArFL1Kt/2
MOWMu2X9AGT/KNV0llM90fweESaWMfZmQO33/XQbYCEDX8IjnufIbhBzPTwlg4LppaBabiO19ldq
34pwzABMrxWId8m/92HU24JCqYZ53yGQtfHx1nXNEe3jBh1lN0r1/ehiIXQ7CiPb6z7mlvHDCn39
FyS6ni2TXP9kZbyZYPuCb5MGdYWv9nLdvmnAlRv+On85VL4GS7fX8+uVLfIW4ZEahQxvFVOUNNq8
Y0WIm+M/xe4N0uFuwdIWShzz3VrLtpc7XQCHV2jyuROsbTkntKWGpekgwwIWCPLHRJvHpcdMUUxl
hhzyv69+7kgjTA8SGRP2U7+wzbbceVmDG3GJ486DRC6DZ2rfYl3KI1FnyjULtdB69z40YV1ynKGT
CsMhWjb10kcnLwAi5qijDd+y1EFrKtB8lRCiZLGFYinVch8rPyc1tBuyiwY7WyWkl3WaDRkIVBH9
9ivnGZaihItUteANAVP60h0aIjzXwvXWq3jr1zvxtKug0tBzRuoqLZv/PDFHZic5/7vZY3Cn8zX4
vzbQ9tDSL1mPsWKKRTErccHO21RoAdeA6lnmHf3NOxEyluszfO7tTw7EC+1xp7uiff/lc+2mcfP0
XDmiFtE6hHqp+Yx4hKw8pCdG8Gxvfqir7dbkawhQqxfB1BybdrdMVyQrk4Jdyxw4i6q8GbRl0zaP
FL2vL+ufdLrXRS9uVqVdrOfTbwOxs1oS2gjZR2DvYInnAYTZFf2/ANnwaDKVvwf4n29jrTP5AYfn
4U4W6rpLV+YxSRyMLW2CiWDQU21r2f2zS6EtaUTwYHlKR2DR2K/oFIC3dT7c+7t7a5UEVC671kGV
/PEyU5FnqHMvcmIXwlxX20K9eLPvfg6MCvIhubRi2WegdnCuF5780ZQ977VZsqjSy0FseZExHmwi
e+LsjZc9+n4Mn8glsPtpVSkelugiydTkHMdRgMabjeR78t/B1NHHZ/rc5TxD7E/y/bGdaJmh5+bu
0Hil7FDtzrIzpnJ1VsImB0T6xgIbxNN/o5AgDCLGKl0BqsU/aUS+bK2bTQBVvKZrKjRGAo+mFKtX
gBDWruEMO+8BTrjQZfsyh6lKTM5DQlvROCuYMtbCm+du2AD68WKvDpi4+LF3I8ad+apV4jVAyMJA
m7fpwJPqgxYIHWKiHHwAfhh1pKtd4MNNgqwa5MI0dN3CyKjNBRi3n7Ney6wzO5lty1vUc/MK6LJS
1qgTTovUq4rXKfssgBHg9Ji1CaHOU0oIkwFscZrMZeHQPyebbf7BdNoa6vPFamBxD1AfWPjyq+nX
BFkmwFS3660paLz3ZwxhXC2l24YNOxEOIBpsupEqgI4ByysvJiJemnu+PKDIzWVGRXv4yO5JDmD+
bUgpdrgZkazTqcCSClv/RMNLoU9UrGezS55eRmGNm6ZQoCoRSNAxK5/nO67m/BxD8vxaEXxiNhF7
asuz5+1lhmFGX2X6ANzh9leevsoDclNlOTlBYehs2ugCAwG5rzQQgWvitfNt90LpDb/nRrYilNlf
opXzPPdFg18aQa9BIUkyoJ9cU5uhxJBQINi2yBhbyxxq+TzBDCKjI0YeVZnplX7DWBpBwP+NGlIw
CpwR9CoDyeOjYapPT8t75tIvQIKDnbLvCL8xtvPHIMQbUm8rAhUT0In+L96m2MhMLcMWTIcJYg/X
ZduNCUkngkZ8y1Wd+EAdGw9YUDBpvUpn4A1F7q6gMtrETw2nGSQtWzH3ZEOfc7/3lNtKSA+XiuBs
C44dfRjlrM0EvwAm3f/IY+/IToS2lu66/8spujQKTBdtvmXGUCaiUmjHHRgb919PiYuvag/r9/IR
RzCRn3AJJsqNH9m1KBpahoWbAd3JBRik94Nif8PwXh/aW/P7liiGv8hoe46Zk1Y3gi1f4y3+JtrZ
x43KUydlrsJOMLNOcfZGujrBNOBwa6cTDKTKAi4ccWmQMgi0XIDmheiadbGePkQTiWPC7Ng0y3ca
fq6UvqnAtkVcW3f5+6Yu0ZrS/pD14YPOn3odmRrY5ZfNGLKs4sYMtPigRM7KzRPutdro5iq88Zcj
DJ9SfvzTGNqQDxUjWmkilbCx6wZQTGFko3r4tb8HuZvZsodcqI6kQGWTDK9aja4yKkT7mE6wOB47
vcInOlvzCmKqpWH9niWGqogJiZJYFnrSZpARu8wHBdno4kJkAxRDWdL+AU7TbFOSUpY6qDdnUtqI
0v7j10raW58VtJTiOIvDmh3hI5XnkjwzLQeJX/wVUbrAMkU+3xsT9aR4QVcuO74MtKayrjbbFwoj
9d5gG02bCNNBbnBBsMOXjlIYoLzIgRqF897ENmEaWtHmG6ykR2UDa3WytMrWN50UXmV7f/2QM5vD
XhY79AcdfT0GxklF7pVOK5F0rwOPMMIIoR01CqUmem+1SFtZ/XHsUx5QdgJgB+D81qQKS4OiZWzl
DA8HYcuoYLaVfwGqbxRv6CcQZFpHDqJrk+OO5qsCgc0ym3JusiReeqM36BDNUQ1JCIVY+mBdHRXl
P38w79AOeN/uy7hdH3ZGnpC9K9RL3VIBOoha7mfg50QSbPhrPaIKW2bTfCsEtJBcV2qH+/44f/JG
a4Nog2TC1dexgK7ukAypAoa+SLBr8f5L0J7zmt2E4TPgOxj0uznGsew9iEEg5ClhcvR4GWWUiU98
X+TR4uO24OAYjQtJISrf2Exb7pSzstZN6K/qj5mCNyILYX2YCXFRZ1IZJka4GTHRO5iDXI29aO1s
qHSzbs6y9XWnKgLGVYzazA65cSmILf+FPAqO3t9QnNoPWXk2EEwl8sNqtD2jMQLB/YS0gHS/FJ8/
7/pdGGOiRniAH2xGFMpG0vQ9a1OKWkVBtzZiwpRMhCf97VbwuiHj6RCD66AK/RQIMapcX7IDn+91
cLwc0OkmWK1UtCSfhSI8Qo1n74wiqu0zwmEjpuVWqWE/pHIOxNRTv8qU2E6aZOz5A30bQ7xvBI4r
zy7XmjMluV/+YS8VhgALcuk9Gy9z3DXZmHupVr/B91LgoFAA+C6nCmu1+oFrNuU8FzLjEl4iOOxH
Q4QxTxhROK4dwMbuUsHEnVGnkxLgcZ7OAUEL10diH/VJsEASMQhaUKlMz8IqFlfyL8tusHXXvJOr
bxvQgtFSqKuaPSi0Ap3xJ33zHG67ExdnVWBA/8fDTFv68zcZ6+strCxD/O4rNiJQZbEfmt7WWTj1
oiyWKBZ85I24ATFGfqAX4qTKc5hX9fty9GrICNp/hxcRv8eUCdTGJIEt6vmvGhb7G3BSvKsUvbA7
k07WgwaahEKRtp0BQG6ykFyJeybo7yss/v0TnObLDWT0Y3Wj5Vi/xWOb+RAMSzNKXDck7xVPoNVn
6BxrmhN3EZoeQMUgoKBrvDHFpaffOTMdZ9ahi+Xd89dnjVL2zl/PBbQvxUTKvmJR+Nwr8Xn77O79
rV/aR97hRPhrndSP6XEwCdDDD+t0sYHaZSOFiYJzDoCSYq15Svgvuydl9Otp0C2c/MZefcL5ltD+
Bm2Dkb+GyGkw4yDJJpNCi8FFKW/STstyy22hWUMvFN5zxEBOUupUYMzLLDJqd3HAxgH0yQ48n5mA
qBLAlkbimsKfirXaT/Wole5Qn/b11fBcrXx0TAkVo1dbuil/IJNb3/Iep0tG5ggbssF8uykgTeu8
HhcYMhX7eCS+7qpKbmz4gX8jqdZby+oWnpVyiDe387ts1lh8VXTSVua+88JhLmcCTh6+ZIW3wIw/
KJYFEmS+16363plvtZlBWsXHrW880Ld0+zYfbEL3Cptxbfal+9b4F2WHADgwsMs+dQRptiiT0rGU
NPjxJwQ1m1WSAcQczi/m/XsReYyX5Hx+UWurzfjkJn6RmFW1JOg1oMkJomTOzxhk6aFbd/7nClVo
ejgb7Ajl3ekV+42L1fd2+QM+7j+ZT+4kuwP2mJJscvVA5Ifd47obk93y3Uzn7Y7jCTdKe/xe4ymd
vDTRWwkeOgov4itoDTJ9dNLrihqs3gKA8rTGJFG7DOXBICXtXLyATrb5cwKd7jsTLhzXhoMTXPov
l/q3VSwp1b4zXki6MSTJwdfhANuuEgeZ24e7mXwpFawQM5GdVmCO2nCeX3jMR0G4gFosDhn5hZMI
EMWVVvCaFWA8OA7SGqZJX0Q/x3xbZMJV2xaRwhC3mSTIqjGOJLEqs2FK9VCbqDd7sNkp9VAhZh18
BsBr47/mo2GnmzYA0LBNIIntQqAkPqAKEeUH+FqxjcecGmOJTzRPUQ1EWf8emH3CScgtMjIHcKIx
tVS94GzoXwKaOzmrEUpP/IYvbCM7y6EH2elPzZB9qH7zUXkOSKyutWpZGXNEPkJRAkvnKWk/+vFk
cOH8u3TvKhKLxG95D9SPLy9qk+iLdZ2vgYmVBLXUiP5npfRhXbnp0+u3moG8fkncIQvaB2sgHmlM
6iH2M00gtuuzKtjdHXivpwhxaflAWoC0/bcbLiRleFNGVRCF74oC9e3t3CoFISw9J/YPaoXPeAa5
wrOo6bQwq0EAln8DXuCG51gqJpiLRozSkJ9naXg/fB3aJWkmxyF/X4qU+zmJn+ySYTlEYybr8vJZ
69RonVuBU+554O8KvfBAlY9L0vMd0xt1SHmeayRnsBCqQmqWk388hQI31+yfB8ucM1YN5tGfGSxu
WlCapBLwbqfA+XAjwSB8DOIOY2N91px3DztXgevW9xnONr/IGySUD7m2emHG30KklQroCFdlntHy
s29FZVwXEqTmZZWyiVJgbboQugbsirUYcH95VDTopQNcLjcgmSM7gqaaU9RN+L3EO4cirsoS4Uxp
VETPDSoHfY1ek7wgCPyTIqtDy+7vhI7mccd2eJ2jBefjgEqg037uuAS7NWqZEsrhEcSN7pK+Pe4N
TUvL8exYncx5/v7FB2KtTqQmkYejo3iJ1BkuYwxOCS8u65g0JZeqAzc06fZTmQ4eFrQiubDX4I9R
MmOs1sn9BYM8PSwgJRN5d5Zz/ZzJwhzoHGnZWJxh5dGOLaYb35BVhjWQvOiPYR5yRBnWMwWZ3h/t
kp82z3OXl9LS6upZsOmhFBUiLm98xJBhISoG9sLwzGonvaAq+w9cEp+NWTrI0/5/rIt1b9QbEifs
ME9NlVOMZ6Yk5sAA6ui6+tG/D08qg6w8VxUNpK9ddnfD+vVHQeqpKsB8QMhV54xb6I+8sBOclAFL
frlBdPvXz4tzHMXKpVEbHpgttLvge+qQEkw008Fx6k7AbSy5ogw9CFhb7gzQbGFFaxP2PcCH5vnJ
RW7F1oObpC2Fz82IAskJhI7OfP4ucVparGDRIgERO/3GLGCKbVP1aDotQud4pc0DrA2+n+LlOJQK
u84i8hfY7Hj3phOuf94jPG8GqYdwNq8We7/5BauvOELLaxX+8Ur27hFulHTsKfPqYWheu6Cm4HYw
gwQ2Ou3j3+Uzf7zD3EpTHwDIGdbsylfu0FJg7aK4zjDYhZBqGnmZU84YP3ovfslu4nY2f+UkiScL
dRPfkmxrJF2XKa3R9FZH92Qavp780t6neaXZzY3YQRFfH5ouWCpuBbk5ZtrOKK0kS2tKUrb2jDl/
zE6vLFovcHXQQT0/cNpuZZj4KNBpyPhbFpptAtdTmSFDUOCOKI2LSklBz2GtGuQJX1mGf2IaakIN
66ez9R4G7nIgm5WCjufAa1Wu6e2pZeH/joItz/V7oYOTatDgSZpY2rvrtxBfAoWt7k+NSKM/pSpn
/qDlXwNH16NfoVL6y5ww417paBtgo4Jso+6su+5qh/eOsePlwre8DWnOLtAa5w7ebieniZgLJj4E
Ldc6F6Vq4mOczzEP7N90m6Qf/qjFhlGP+ZsM8fDfNVMFnLfrymayHkEBnETo6nkqtpyYUVMWgpJ+
C1Rb7ZKD6rQTSkPhBcRRN3bV+detd8Qn1FTxk1Yxq6G955uQtji5UrITeo03Ny0aOudeFsX3mI0+
H7tXOANlhPEbpxuOVoBCodCzR/mbSrmduDEWIZ45wkBPKoa2VXI4GNgAu4DdvL8pVMg5dbesKqH+
ieOHXlAHfBlwD3qX4DU0FqPiilg4Zi5rqWux2r7IH6y7FWoHQowtuWgWuaTDeL3L++ckOEhEBBLz
qCr1BD0yyiMMYdFvZDzWdxRhNGiwGhWz29TDPLfcnrvID0jw5d/fDw7YaFA4H4cRyIZoxiWgZO2D
Bo6Cvs3GwzG5fOGKSn14sjEUr5w+ZqL77O/xzaxC2sEBGXfQe63DHuvbsy6rXPjpoqpSPNuSLQvm
nBHaSof3/A3WxuO3pHcSJ+hVoJumlBpWnMe3KkX3Uo7Rbi6vM+ULEwtKF0PF/LFYdHlO51B5hhYN
4bQ/lprxtRRm6dNYKFA/D8kVarrz6MWecpO0y4ajsahii+l/DAiSBf+yB+ZLCozyzZ2+R8BLoOBq
lytQYOP5LhK5QqJ1mCcZJPPe04NIORuK7S4vNj+heShMGAaOXLK1qM/lLOXIjhed9rqpmzdSYX/b
p30anJt5nf90tBbwX9E5RkmYx8UBbgGw91zf8Uha/1q2/M/TexJ3SwHALAEjzOU7T0GfdUZMh18k
AMgiFrp7oMnsuvhHNw8Rv0R4KsS58NeI8J58TME+zWFJ52NH+W+cXlO7FtbjEpWfD19jCUXDi+f1
mZ62HMSl5HfnIrlkY3ang2J/GutZF9VJ074zkXPonWkmYEGtRl7hfdyZXMWlXnjFNDuImTV62N83
gfQgAXVF3kHovwxi9yGMvqwXDaXyOmFQBXqAbStK9jqzj0o8B+qzhqYmvIzXcXnLNFY5QJ7ppyVE
9S3hHUk7zai9ipIcTj1ZCPl4AFvZq3S+qCkKsRQKOj0lAusNghjpdeK37puKvgk+7q5rXpKTK3//
2pze9L0ZyuTTL15TbFqJhABC/+NboV6uiQro//6Gf43U8MVt2KU76zjbXR4ulybj4dFE2Xn9KWdw
cVXTtWX5Bd1yPrhzZRoFIHv+prXnEyJupfqpaAjLyxiPo7eShxvXP4mGhGmTg6gAFKlBl+wQ4uwT
k143IpURe/CyTOPvWAzZGJbSNabOL3oVAlVCjpG63sihWnFatMwI9no6TlS4tTGWMjqqMaQUkjDz
zKyWoOv53/aiczUICGtsUnAa4BKyZJ41gls7jph+g+l1w79wG9Bl9uleY0rimIFIflNmwGAeJS2a
1Iib5yPz1p8pPCXiC1LMS8Z1a2zj2J6XfYd4D8R8jAAjw8rFG0rmWwtiIkz6ABC8yR5cebv7IMD/
VDZ2JhyBXTU1CuRFlQ934cbzmEAsaiSqTHRpWcDTHYQCPd+Yioux6F4H9unSaPvO+9aTVHZwvk1Q
vEG0A9kXAfSKFbVjWR+5azfd8Xbk3ESl9pxQ6eNU6sPMFHHPAgxJrYNzBu0Ayt+JyJ3EpLsVMrWs
pIzp4uIYR+BJTHj9tkBAJm9DEx3HNInKnHf+i56pp47ueUX+0erMNxAj5LNpkBBySuMhXaVedGgK
9r0w/nblZ8IQtdHJrksyqKDIyVpFsfNCJw+VWdJ5Iw62QHlRPxPRKKRYBkXK5jflAQDBriLL5WO7
G4y+nbPNpx8RFB9C1pM266QGjoBwF36PMqKQzC3mfFvjAwXUQGVYJGefhvy2WMPeLnzfwmuCOCBL
5pXtvvGnacPf0r9rVqh1Pegthmi7KiacamSAax6GwZrNKNzFE/SVPpReFrX4A+qAXA1gwN4bIyZf
+3y0I5wqilb6ElTW1ZFXxcJEsjSaPw1dClfwCmsDx5LTE9iLi+N1NeEj4S51rt3L2xYVywGnF/3A
a/U2vzFE6A9MXMMlz6oMZXluVhYLMDqaJtXiTJBp7XZkmUhWzrDaPrQARlEjG9Ww8XhoHthhqGIN
D26yUybwIiXOlRhVcZP7vB4kAFGx4k+QgWHAv2VVtscuLftbmfY7kxs7ox+4sSCP2o36k3iWiOzs
SVH0LZkGISXSs9Pxdmj1JZzgsKiTapPLPRK0h9+58OC4ipzdXBPgt1hkFK/1AjPBRuaebTkaRc81
Qd1VHlFo8IKgszMSlk3OOSPP3rz8fmjuminzBiI6jvxiwRrSHibHClCWfgznXf3kFbs+6/mnDahS
BCBetVLOeoWnwLKHp89rUC7Bx5zMwG2o3zNYaWfwJZL4HhpXRrorM2psyQpGlQ/8tWvV0tdpVLBv
zJx971SKM2COJc9u2oo1ZNf4mo0rWDwsr32jZ/q9ydkA/cNIQYDJZArqxQETqB763pEnmDpmN3Z+
M50jHdeojZBX+37d5vXk+uuHYADxt/XqccvXCc1vyrStumBS10fZzreSF/BsJOU3T3G2NvVKPi+C
6n2i2OxmBSUmTZ231LSie4+PJHSEKEi3ZAEeKcr3YZ+AbLu1fN6cMcrNyTaS1GpUQ7wN85RocZ2Q
KVrIWMt8ORQ1kIEDnpoxwj3ACTYI0TdkP/iGUjrpzIiPraNUd+sMBBb8U/JUL0LmB2pYyIAq2sUG
GCxCkrB5Od7mVRd73hm6hnQbwjNi9ldG8r4JoYeeAazBTPLZIj0bhtTJXuBpcDdiPkyF3VSfYlLX
LqEzTPK4vGkH+iPWJt1s8X4CcRxiD82FwCH67u3rhru3HToL2XVnKehR1iCAMCKIDdXIj433AUZJ
mu8OAAxAc9vU8+84Gq1+90hKwrWneKrT0R1METjDXNz0WqwzBBTYlXUqbNQwsSDMExVyIPr5xaIN
jhiTLfgwEATAZjDpctWPvtHsE2XjcpOOoJYFUDSL9FEIToFgaHavz2RwA2YBq3j6mZgb5D0UNRu7
7lWca/WyegThPTNd7UA9w71papSKOrxQKSsajSLHHvYbdKCPaaxYmS8rvoD8IX4E3z68+4jXTC98
lVWbD+wG9lAKBinmQMEE6kIpl/GE9F2BwKbtagAq6nl+BWlkQEnKvc1cMQeQ5oI0mrAL0VhbxxGd
TeZqHQ1VGIO/WvJIrvGmtL4eDUsyJ5P3/FI/J45uicS5ejnjki25e5ATk4a7kcl4lQRoH4zjP79t
uFxQUwsAEQ1/konNrlgCOd6gbVuzMxYeKxkWXYnv8MYXDcLRNqZMId8NR1ibuxHxsdmsryL9n5pe
ChG/eO0005pLxm8c5bZfZnr0SdQJzh68hTucPz1dhGxT+uTr7LN7c5VUw+gLsoNmgQLd+XtkUpfm
ifUYUA6liFiGn3Z1GQxfl/TMN2muCe7Q7Qgz9n3jHCg683vizOzCZbliFHicVMY6am6NxGFbBbLZ
xHFc7BwAOCXKJhOC/OhODG9x1tvAzVwUiySr9Tt4VcKlUsDsDvNRjVO/KAq9eAW8Zs56ostLLpW5
U9kF4Y+5otHap45SUzJOBbyq6J9WsuLXAJQjKVxrZiHNp0vkcI1sBQpGiS3wz8j4lhKyek0lseRY
vf4ABRzipMIfJ+hN8zHTHFB+0w7N6QXACNrzMLTyOXPIYqx0ufkCb6TjsCo/MW4K8b05t9uqkV8i
GgsgYkf5XB5kLLVBSVVF5mcO3jZZB6uOOSF2AZJKcz3gYBNHaakK8ttTkcW/jdRGy/W1vsSFMMDM
jUXRU7xBDtYBiYZX2cdzkPvucggnmIIZDL3dy2byXks/DAYG5tVm8oMuKG1BJ5uUysuV3rhySqLe
OCCZGlI4htSmU3/qXYxZuMzZlqtsVR5VKrLMSXmI+yUNRZ41UcZQOZx4QsmsFBCZkSIJVNGX+bk5
80ByL4lkROKToCzFNcbZAkx6YMo8cX+TEeCabO4NnSu7a1uKjTH4DYzMTlIJ6f/wKJn27OrO3VIL
714i4y58T+sA771hoNor9ApzVZK1HyQ5XBB9jz8AYneuw5sBHi5fj+Vi16NVIR9aWeh/vOjN8PoB
wUMdv6exBKrxoh1si++LrdIcuXiepX3KeFnBlXeEpvqTqUbHrC/yhDGpagP1kR8QowoiSSLtaC9b
vhD+99/gUIsQWG/Pru3vm/w0QTynG0yp9cblnEVpFTyVPSFNiQm591VCUV4azurMxZfIy6r3W8Qm
GOmbY6UfXMyMNd3jrS1x/LqzwG9UsNBnAeOIU97H/d1cHVFIbnqHpaM3Kjs2kUfhLYDyl0eslb4S
8kHprxjoHd0CnfLMj958PokZ9ulCd2QDBms37vk6hT1hdHb+tDtRngtpfaWkd4RlD5T2VZ9IsZBp
+hug7BBKvyY39lRnOCz2dfyVdhW1mtfDPxi3jRwrrwlebvAGe9eTU8sd/73SJ8UEvXIiPLtAIDVE
8SDvGUZ24+SjgUf34N2Rm5H11Sb/KiC+SkQIy8T4OhqBLH/uwouU+7e1tPPIMcnWJ9ZDRm0beiY9
lNYWvxKiyX53i96gR5OqWXOp3Y2sdH2OgURO4CZ3NMgv0Ds4g5uxF93zzsyPQBN9m6KQlqDNC5mi
nh2F3my8SuIbH6F5BxMPyOuvpSWLboY1jHWbtse7VgZm8BvyFUZPwpP3iEMBXIFxQpsfaUV5WGuN
W4R3Vdl0nGK6EGql7iESHucPQJRltlU6rNDEzk2/LY0I0qEZFkQpbxqnnntpYYPKmuB+gHSo7+xC
q0TGSFlRKt4QSFVmR6vK5x6FHSkX6lcZ6rYabU3GelM+583zFWkkfHzkvfd4poyK5JJh4ceNsH3G
qBCY73SCBjv+2meqg8fmCN2HWy9O8GV80/lDMwpVFO7HlpQadDG1tDdP83mpoxvc75MQzOkWyzwd
vEvBnlZ8CWbCXt5dFMxT+pmqH0oAuz7TiffR/KEK6ZiWgGGsHp34LpFwkKHAAC8CIOVBYAVebrUw
BDEMJYImCOVCUiVAvsV7w39C4Vq+jifTdYpfWrCAaVB3qoJJ+4UPGq5TpCcytCPFerwhARP2DE9/
Uylx9oyIgS7yOwipXN1esukPI8oH/ul9LkEukdzNSsrUguddUs/3KT/Py7C+J/UfQ13klMMdKDNO
gqQgS32nPlurD6U4n9167L37Dx7ud83EPif/ASHs3J3+cqtZu6OstV1dnvI5fyI0Cy145ecUr7vu
TdA3gvLCtgKQqNvse+zguyJlennnvFCLwew00kYouZAPRmNMavpfNsvSQiRM8k1qvMbCUgcOtUnq
aRMFTRj3INEbI+JftR5SDglNILM43RAg32gt4aIC2LyFH3NVCM1376ZrX2Q+2lTMmTrQyqrYEA4Z
oVFt3kvuZP3kB9FlpU5pkfNUicS3fJS7GELmeWK3pkj85NRpLbhlN8Wf83mRDYwBCOSYZVRQ0Ok1
L5sB2q62dJqvmCskeoVNqBkqdiX+7Wp5tJyeYA8lsx3ojZv54qzX5OdWdhs5/UhinsZQtxI5Ek1a
CO+itM8331Zyk/z2oqP0X9TH+ivBmw8a0KTlY/Y/GLwUhNIhI/PFz/2YlI/hg7hiTtCypyy4upYL
JaivYBZCZG/9m46/PaG3QgkQhFVEaWZB+GKBlTI3HMFNan1o5qnZDu/uDw9lftTXSl2xac46Jca7
17Lj++VYivs8c8SHlEzGFT0n2IpVBCX/nipWswg8OSc/++7inJ07YYBUZF6WQKJ5Qf5dMWcIEVyC
/0Gu1cs90R0jje3sfaqo28pgeS3f9Ypql9jyv1BmiH8Vui9TD9mI0vJnEuaDFoXqtaxlT6P9Fafk
5Rmks6tDtlmOdF1oh1C6urevqDStV55fdLacgW9aKp6NybmgwQjroYrenWXqLHKtkGPAPBPK071s
EHEheAy3VCD9aTcspv5PCcKvjmlap0YkSoM1KlMQ6LToXjn6hzE8/i3zY682m3DuCqrtYHZUheoG
7uXDLeShUJ6PVGtx4S18HUov8mUZNSTqKawy/X86uda7QIJOsjSpQpOuhkuDhgXHrl7515KYdvLL
NDCkvx9UkSp41m3Qu+y3i8kzekpimLuHclqU0gRkI4KStGLRlQf7TBJKbqc/p0AvKBkKI/7VthBc
F8Vs3bP0B6F/Sv/sbLh6330X59lNAsS8WA2SJe8K5HYv/9ryDheRqUpxzsCPb9te+vrfkETs/6Tt
NXmuUjLT2L1IEYpf+74zfY8Jt9E+sizsEBMqhLAmSKtE9SAEQ/HqYYBaXpZjy2VDL2h747mbap7A
TP85Z35X3nAs73KzUthwSvLR21R6jZX8b0Jp0MNbdelxkUICXUPqejM2CRKBTZQgC/4quTeU2k4c
shav+JN+4oEdmldAxW3dt8CPgAkzRNNrNsqhpc4PhNhf2vlmflJJC4LrCuTlQhhb4rmafGl8D+FY
85YxRl2eyi7Op23vfbZJR088PzoPmxSRLZGMsG8vhzO01WeeEKePTiKGqZ9Xna3Yi1Lnc/fe0Zp3
8a+hqYMZ6M3cKq0Yo/rsgkDhkkyos4d/JqZ1WmOsW8PiSmA2HZuWJj4nVEJ6HYdceeY9Ub3bta5s
mnWXOg0HcDYf1s6joYsGMLR+7CLF80P4w/40uNfImZWZqs5Moy7q83FS4ws2PPkkCTq+gS7+Q+Fz
p9Xy+eR0+SKf0SBvwEboRNNGgbJYwLlXEoyJ4TdkzdT1jJRKu94J8TVmemtmARNtE6pNOgQtYRCy
roC3+pbMunbCiMgcOU3L5D7faUFqHdg9d9rWJ+oVJCGWclPlNw8ocyo1Z2a+AfyvMAK8MwNw0QsD
FFD8kc9ozE64ath/AisJ9trL6DzvHOjbtI7h+VzCCNr9oufVw2CeTvnesqop4Grb0BRfr4jgF6bu
X9Xo8icE0sthdol0ZCaUS5Zm4cX4aOcPBJM1bNtxXMxroT7Z91Pwiy6Hhl4XBbsI8Zq6PKnnkfhk
g6pqdQiWZt7hs8iRfXoEa9cFv3dH9gffAXrwcodxB016MIjZ6QN5HS9myNFy7DPpW3gqpSxoTdoz
Dwi7OpNY+NcwNx0Dv1s8c/oLKAQ28LlwxqwWbcIqefhcI5JoXAamgqK0HLFdC/u4TvAHZYdOc2t8
MxEP72LWdGN4psoThN2F8adBet61C7knyFBJZ97pdCK/kLjAC4EvAifG0sLkODChiChkL/iZJpna
zh12dIRZAtmptAfoqxVkcbSB03RwcaxHSNMR9pXZ8lZqe6mSCioTryZV6q823CEdGEfJZu/nieSI
YdZuj9lknX4lFN0c2MVjyhu34SlHi304ZtGz0ivKV6Vn53jr2KOZvR1Fk0chTolkdXKBG3bO/les
wN1sizrT1ler5n8v58Jtq4ju0TaIxBYT/UEoGH8ETTuKLg/oRIwR6iBDGAu5dyizjt5RfoodTuMd
hc+osJQtqZa9KVtLnCCKeDMBOBqHuiy/GHznxjPl4ikm2iDU8bvgj2gAfB/QuejWpvRJLT5D9CBL
iLgJz3/PI1M2PtzQ71aJGj/ivGDZWKe+QJp4gttIIGqjfFEpBMwlC8Ek30doocB0fbAwuyociQGB
DCcLD2Is9xTRDhcSjuVtVrtC35Kwwm7s6/r7EltzBRq+QDztSdzr9qpfIGPZf4ojYIbZa/JiqTY5
akB8HqYZqIDMNwpEMT6imY6kADPvvFYrzeKM4cxNopTI7tSIPqj7fQS1vYI3dLqfO7+Zkwd2D7D9
hXL7ISh2tkT/4RyRmTrRA/ULRNRSqasgxfAPA2KNftKI1a4JG9pKqLhE5ASzomT5ttFUBA0trQx7
TLAsZEqLP1vwUOC5iHFR1MAKQqtnHHEy8q/E+mV0zHMwaTiMqEywaUSI3Vg2ZgQTfLfaJeqegwIZ
xdxQiDO73g9qTPpnQqXZt3+dfTbNJZ+l7OGDAlxTT8QRnAxcF/laGECI0xc2OXL2NRIDH43O6kDZ
20FLXuTPyvEHejjPEELFCjbtxNScwsyQL+tJcUwPNoC8G4Q59hsuqnzJBu+WVHe6pnMgd0u57rCF
d7iLYo44/tZpFNeE3VesiEKbjGEpohuzxqO7Jvhr2eba1EkgBLvRZ+ns4OstyHHgXq1XHVs7JKtw
rdXvgTW9kvI81wjLu4ttKoVoIOzCxXXz5nNBOXBvdnUGsP5RsBd7TWt3d2dL+YMLLnXJ065EBlOE
IRigiJnsYj4lwNuerYpjbtcqYX4uO1LML2xc97JPIVxSXxo3LASYDdAof6lZry3MwUEwUZKrIB1Z
afgeI3AVzCkxgMR6fr8zIIf4WQjIiu2K4y8OO+b+yQLq09lQ2GCDmrTn0uX5lLnZWbgGFWDTidH1
oPL4rcKPzHVs/m7ap6cEdFzf+bxVosF3h6pu4JKn7O+ZbSnSAyZlYYYz0cM75c49Sn947Sfc8tLP
HW2LabcYw7LxkMEgIJroNNSw1CH4WXR1zK92Mf11HDxA39iYiTMTU5LGcsx+Vvt0kRkYdKIsv2eM
PpmUnEnmnGcAKLvFcE2Y80D6DstMzG6LVGIj1FHrYyDdvnU3FqRp78rwu/QO7dTYLqgkx/KMfaas
cFOIJl7gxbed7CKevJcaYCSB3IQ89nFBdUcRoNF7xp3ao10/VDs9eUT1Ua4USXd8mQqVAtuuun4f
33Cu3e/SJFa+EwlysXpEAWJ1gG1AYtD3dmKo3P4+fn8JjQj6/32i/e7FHWCszmRzp+FYWjHY9jv3
41NW9/pXNFV9j0d7yptwhCbljiewOeDxXJdeRFc+sH6UZyvU9soCEUloIV4P2Wns5Fe9e1lBgw2e
0E34FZovepFXykBnuTfUcsJV/jlxNEUD9O5oUBUfiw7moztEK3suO1JNAudKYvbhH+M6fuk/kl8H
db30N58TO9H25vKUiEJFo5j8MYbwIUPAmR5VTe1CbWbJDwpuzQ1qH/x0TpN3otzrZI3TA5SuUAHA
9wZiw185oHv8GfEuirQQNWJ0GjYMS6gVhxMjkXED/0c99yT/cXbj+rACqg1YS30XGDn0cxuEVcEB
SmC/7PwucmUqox0F7d3VYICoIrZFncgsua0gynsXEXPbOc6yBQxSJUAJ/yugh9AwkxgDmieNA21d
TQg+ZiGVJmNPsLPV4xfTYgzc2/Sae8onJvM0jnMYinoIKrFwiLHN8jVx9EhNpwwKMXYTPL0uXaLz
eGxeEV3TDXWD0ontKtOw72OBq+yh+hYfGSiGvsEBGaqykNqocwUYOT1vEs9iQ8yc9aJtzJ8OT1lq
hT6kLx5FnNN55twSw7GPFx3oRSgpjMee3DzRiB6Tt+0dV1ZcGplS4oFDG8wSazWN8Wf9dgRobNZo
FKfeW3bNFJkuOnKI+hqemKamEPH/FdKdzPEiH5oeOWp7e2QNg3ty5dITfPXL+dBllHwrC7eP8AMy
erifKAnf9MGzlu5Y1jVlWEciPD6/RcrUvhBeH1HDtq4tUcahhC0QFniuuV6VCNFJyzmHerdZ6L1v
7Y5y4mFfhSp1HzKRX9WYmLCcgKblYmQAP061I6Yxpe46EhZPncYCOg9Wm1tcgC8qtf1POdndrPwg
jCq9FlQYkru2hSftb7pBixFF9ZtEwv/V9G02jEvlxfa3NFRhjgokhiMBfbynjOLrYEV/sjymabGT
buHF1yr7DO5xIeLTqnLIN3J8CE6UyMSz2ayptgZ5Rnmtll6wFIEEoR5+aCYzv2b27o6GwnAeZtyS
JN05f7TveUgCzOBBsF033RFsFiqKg+vcl3bKfCG4vM1Qgveal9Z9T1HBbjXCRsOfW2zAie6PYgzv
3ShnGcEa3cmRIfZjC8bwESVCELfPh6yZYpZmEIMhArPHDJU2pXHWeHdJeUGJ+e+KM0BTadl9kX+x
qDQMsBWi2++AalfNppZkMygrvOJpgH3aV1H4pRA6U4glxzTSxPj58H4inUAajcrBnyacwpRrQ48O
stJmYA7rj/Uk2umLBhHEdzw/ce8CgTg1DZOTHFm2cRBM4JuZmDqoARnlYsiQwXrlrqF/+YKv1h1x
iCksdwndsHjU6RySp1GJRqVuWaUdNiOiK6Dfbd7MXOdkGS7w610saApkDTmvYAlARQJRfmebk/6Y
B4E8pS9KfN5nREEKz6PQLqCaepqK4w5xSOriY0yNBOHxi6cctATK9/MC554YS8L26VKEBKXpI74l
KfIuFyL/x8snWnM1dTdfDww9dbE9Xm4syYIuaeP9MKFJSm2CskwgmjQTlu59GhAM3Ivqz81OaRRz
GcRxBCJbhaFFTWoqur2zgq71Of9mI1KyF7U/Gebd6cYhQCzkyay8eoBr94dYXq10cELhhNSEQwMi
TmdZSxTkXLNlBAhdmPqct/tLuxdtGq72VQ5AC7tIj3sf+ynJCc/F+dhzjNlt67W3u8xRXTYvrJvg
K7dsEpR9idXC9/ZXKz2dfMBfBAJNfGapDu1Q2t5NyRFRXrxUEJC1N2IDHICrKYoM4wNZYckg2r7f
Y/HDkCo2AugsP7dHh/fg0tdLKJi+EesSvIuuEnPYZbfGW957j1rqlnbTV6NcSPC5ivyaehfirka9
Tmm//RO/CCBv4zqVaj5bRW2jrN+55lBf92Z7rsrAtp/MbkosWMl/MPrHwdHGq14rCNtx/W3QjVLG
AynAItSHNvq1qIWyqO3bmR57r0rrhumZ+1HmItaw5z4Bd3On7dvhMytR/G8smv0McLjyk0s4QKuZ
xC5bEp7IrxZZRPB/mBRcltYFFzm8ifwleMmj5WXsyXcJ3PzyUfxM6LuAneD6QWrx1b7rfgHaIr/S
YmnvAWuGVXjafOkb1IpwpYv6r7G3UtboTzO6Wx0+zPq5QpJa2rRmDEdVVVYg6XD57E6nt6oRCAwO
WEFgnsS6zFN1yIXgNR+JXFkfrI6cSYqfyf20dDFN66ARpRypBdHPQrBR3aKmsMo8+RRvkbaFHsp+
NypjQKoUFAGu0Fn4wlMcpRq8Vkp8cWee4q+9nFdHS9HFz2Z3cqrsKF/JdXTgE5yO2wjWiR7Vi/OS
gvkH4SSpGy0w2jPudzHHcnWHViDsqFfLDJPRd+IdJQA2kzQ2UhLN6cVg1Ie8EdGZEBOoJetdZhpF
S9TvCew2pp5l2wDDILRunHSz/7ujH4dyqLmUymbmnKUcWDhznVzjX3uVu51LywC2hDAEzvi7C/1q
daP7V8y8DGNBDNaQ0Obx7sJzHoGFn+k0YEfWmAef3cxcw+XPv3f6QRpLTZWn1tmnJEpD7Ojm16IU
gqkzn6UQVWD2bUd/R7MM8KjD88WUaMNEK3Y8z192EFwViidFnUAnZfollobxld+QfuFCemWHhfq/
xE1r4iK1sqjAMu3auKqRxKemzfdtIuysaOGjpsJ6qz4KRGV2bkiQyaCXmtnIdhwKWBUS1xpz2dRX
vqrGdr8R3oiuMgr1knAd0t5M86hCwWwGHh1oWULKDlmj2Aq8dsNE6V1OiEIoJPC//2XcqUsZsubO
uqiUctuvKjYru0GHzww/9WUeRObfP3u4yn0Ia5gKQi33w9+fpBtMN/goEmqF/bbqY5RoOXt6FUzT
bdnmwtu34vWyekKHUcs73JwlWY8wMAJ8qU0PwK3TrSsV3pCDYoebqCdOtnk9slwFS9amHgw1cHxG
r45nyjT6HGXgzjPw/twnI4LH+Pmqju5q48+4gsPiP8/fRhgb9bIaT4T5cioW1yQx0YCRLKrWrOs/
E8cDKoyNlpQIe03FMrc1VTQzd2Vdc1vb8bZfGsrusArGpHWmLOPPoXCcY0gLoU4WOVAeyhhP7ehJ
ZV166TLlWtzEcUKIzknr1yNlNWUVdpsyrCLmZAj8Ef5V0y7bfpNoIiG9g8jTOukgytamNeg1BfZo
ahIylUTTMlEE8rQzOZhbj8m38GaYg4+aU6E8V1SfBg7zlwwkPz6zhEuAjI+1JE458x1OoHXomazw
zOFIHWQvh8PNtnuLH1Wq+EpcWi69/AIs4D0Mslv+GvfbR7ppSC9nBUHLQePZrJwfP6rvG71KQSw7
+eGnJQPS/1GYx+AmoRsg8pGvFsRjqEF01Hru6demZSsBzJLEaPaBwwZNGh28r+wztQN/xAbnMvZo
kYNkf68LInzr/jOhHHSSiyzXfj2IF5Ki6idKqehC1VD6cdoSq5pwPKNkFPvRTXwzF6bqML9YSOdN
KKj55bfv94rouE8UztYVZpRqloxaAGP5+Bhb6AIO9bGZMqSyio203WMuzclsa5PCbkgwJ6JV3VCB
SVWzRqL9RC88gC01TEca8I2dSRHPfnO2fB10s/ErlkrPxoVX68JWHB3tFbsmX8SXyiRXyfPTcrJ5
mohc/0OMiT85AE94eoKA7Ny9NTX4VHPN+FGaYcAyx12fqSIVuZaTbunGn9H0bBCbtN09XNMtBdoz
6icFFRu2VbjGIV8Wgv/eJ+cPBcC77SfXLo3cLz2NjCiGyQF5SHvVp9HiXuodk5QaRSCr0Ke1r2+v
6pnULldOZULB+5D8Qfg7o4h0OtcL/BNxK+Z7QVEnOkm3mv5XFL1nFW3mjdYM728yyJv6jonEkAi6
A4TJayjmGGd7r8ePDA9f+QBF5ZR23UNz1pqAbV91RAUr0OgUx3zx646voabAIvC9TpZrgUUpWeJH
AEwtz4bO5pv2cW8Bxz8vbUK6rpHxTIBXfCchcosZL0gQChoybFThNrYd2V2OCn9JjJbSySRote2r
npBU6P8Paafvan2PWTAn6t4NP0SRjpNm358ieeky7ozEpS7XYUVupJGf3p9Y8Q2wqkRcvO+zdk0p
fV5JbLwFtPbARIOiTTohA99RiBDE2Q4w3Ei9vy4zXPT5gglTC30Tm7+nePSmV6NsLXT8VwC/vkXH
6lao30MDbkvnrU27x7F//GR3QM5WsVYX1SlHgAC9WTZ+S6PJOMn+qCRyUm+eRCB2PMmQh8ohHVJz
RxXh/ZIuQVNdnxdDY5I+kB/eSizeYXGhoDpiMFtPPGMr2tO4cz5IvuNXZnZ4IfwLGZwzvJ2MgA4s
ouYNiTVdLmL+FU20DrHvMVakxIQ4VM0Dmrw0wUbiiZ3YSc3aUPw9dQZFVJjVC+Pw1mDT+9et9A7H
Qjo5jaMQ7lmpQfUoVZxPF4qCpgo6jbipuIbrawjF3dYsxK6XzX3JMcC+lx32EdYjUUnxhWXiEPtX
6/PUN9NXV/K5xvfBuCEsdLZeOtmS+oVs3P7nkVYF0bIY3dYf93TCdlb3ecE09nh4ceBoOrRiz2WK
NWsbC8p1Axh0AqVnl34G5GrTqjzwpiIQ67iscbY7vwNAfjRWoOjYa5fQZIrFpyHiIQrE1J9XAFr9
KSao+Q8hxVFFuZwSVyoXvW9NgrBKLQkSki8FIdjaf0QEhtOCwG15VCHBPw/u0h/ZG9t/+iIQ4dP1
V+bTp20AC3IC8lwV5Ft01IhAGV+GxsiyoYHoeDsiAXqZEH83LEO18285j76z05/QxNmKae5wy+a7
daq0iBpdmm2RBsJhfxc8ET10l8bqaZL42tUMFDoErfChpWyh0dOjiM5vtg4kZZjwlaw150Lc84Zy
SRJNHPuTB4x/arSGZhV9O5V3b+9fyY4ZT+80finX6cWTuAROWG4YnZmJI+LEgDvJsI2w9k0kMPs9
19VnNeMMb3zSVoH7s7BITBR1Pnyw6SGlhmnfS2tmndd6MPUbXi4Xcura1Nsp+Ouau0Cy3HlNDSvR
uf8O7UaEwKYwiLtlwRb20FLCmNxKx0d37lGm62an2ZWSqgZYLWAzGImzIJ6lJV9iUmRGzjp9jaHG
JTaJbQQvRfekPgFk9U1kB/DGDP97gNJhUUHxW1No8hBSqeSRq4DxlRMCjRQoKJE6Qhn02DfcNiIx
NdhYIQyNZr7COgxnPT3eJ2Af+fMh1+4vCSPTjgOVdFHGCpSr40L1JSjdzX1BtUZenEbkpT1KfCd7
+loeZbKnQcBatBMeWZXUiFx3S7/nonrVGYNmI1sh9YOOfBnAuCaxYFZtSLEpXjHZ5Xad2LJ1YawH
GvN9SipcUQ+QHQoaZ2Vlj7UWBa2TX3KTCXiKQ3D2fmR+Q2/Mb55S+llhwsSsiZOnN822WFBdxvVf
HWMQcD/y5d7kfq9QF/mGD1xw//pjfwieK2l6fP+Y6JS6z+1tLfOs34SJ+kQStnhGYOHKIRGdMtFK
8cWnthXy5Ff1WAQPLxAu8dkOKDNMGNXTY4XPztN5z8G8FegM3hulPx6+evvBawxc64NIYeKo3dqa
D/zsVZqcq7+XFPCuo5gsj+tNAuUxVzxWTieq2cNqT7FxFm9UpGnz1hTtLRJvw3pKqor74mLjkaqH
fX9illKF8XmimrRv2LBVjjPNwnmnzS2wlF8B01sdyRxyMyIMtdVWZkv/dVxy+B0hkcQj18h0ehup
3PGPFgYPZIjNsBOCRvjVlHmsy4j4l5fALQ1VydIsngnJobIGIU/dV1ceDGjmmtBNJH8lnsIEUOFi
KJ0Z03JqPyY2r/WlBeyQADVaYMMNi7ZkaBfWLi6PIe+zIXs10XZsEqr9RUxerEMFqkOgC+hrrgxe
ZVNdirBixejW9aNo4UD6+dvA+lYAo6z9mjTx8HrQhkeZLpvrIXaWiYUASb6au0dvD70c3o2bz5cS
6cUGZ2af2d6VVadtrEmFmk2dz7x4AT6raPnfj8KHYQNfgccCuKszNWz2svWkHTtjCFsYxMAaxeBF
7DZ45RuDkSwSh3+WNXz8QVfrVl+uIOUn1MyHkY7GUOoFDkZwnoeGfa8pfwl5NFfTYA1S9b8hz78o
bNFOt5FqBVkTBA7t5GuBT172QM7KVgDt0O/wb3c85m/oGK059sfZznJ3VF87EBTTcX3UAxexWZoa
g8Et9BSI8xV618C2cGCTUvsy9kcb8YF9jWBfilBny9GuM4aXUbggoc2VIyP9Mc3+s4RBU0IXBWnN
D+3dS/qpKKqsjzk6w32RcAvgvWrtTue3Agd38yQXMfyKmuzjKMQC4Q4wUOQTP3jRCHokqYmBulNr
e9L7Xs4BdXdIOsoL7V8XVFXMeQEU6XBFG1qAIAPJW0uUkxQHIMDIcf9E0yQglz1JvPuMoSpZJl0J
nxCxxfJ9wcqjV8HlvdLb4z7qrJc0NIlMsMVhUE6NHK3GaRvnDXcbkSdWk9txwhlWHYCcK/Zgtvyu
AUYo25+pvwJRnZ+5Btk2/aoSMsREpSs5dhQ/j2zJJG0hBB0GGt52Y8ni8WpvZJbktF47grvj4NS2
06Xr+vKdMM2rBuLah94+yFA9dT2CHTcSnGFYqWnNsobd7fH1byFW2fDAs21sqq0vuICF29aVOUzp
cLvsR7+C0z8zdXQS/tI4Wcl4E8mtMrassyoMvmIennI/jctH5LphuMPgP/3iW5yi9EcgX6K3XIB9
6eVhUrwQkTK2JXnnRxalzKOUk8dsFtG6PA7kK7w6G9mLKWQ9oN40H1juIIWXDcP4m6byMTnObuaP
BJWsYoqsz5OatWOqc+geysKaKZ84iX0mhnerXcqbOieLG9cX1VLCd1A/h1f2nmM+vKZxru6+sa24
XW0tRO2Fic6FTKFfC0Aur4nxubXkvCzcuyYPbVjI6A4EHo2m+kgTCiRCu7FQDKq2IRsH4Z1vm16s
WuU6hh/3faBODYJKwq85PreOgecV00eFq0Hl76DeOAZblDAIKW38TIIWCZuHj9GSFYDiV3X1J2PD
xVtpzNJOCaIx6/81Kc81PYC57icELSMZa5XAFjnfFMRU/q+x9NOInwwpeIo6Zl/KjAh+w4X0AGU1
BM6l7FTYY6JOYz6158QwC/az8jv2QeiOWXfr35f5F6WbD7vNKxY2KxvlCS3ZMkie7nFbdNAkant5
dHmhBXFvdlf29F91k4Y8lwtlEwjE64henL3cXAGLO2oBNlK3mMtrv0VA5aT7GAhU/WCVhW5D39pF
P7E4Yhz9g/Ys3OTe6U4jwdBIHBVlg7z88abntKsM0IiEnXap9BfglD/TuDGycf0E1ifBrMbD7B3S
FcXOdzk18j3p7vjlx555D11ZQVlHI3Kz6B9+zPDVAUv5saiEQmDOZ94kSOlnYl6z08U7o7XIIFx1
H+/SislFb52C/akMtZqK1EcQh5lLvg9nXW9syQEm8FGmmOBw6GmtQYyrj8lUS9f4j0PT5OZudphJ
awFU7pgcVPOoht8J5sZhr1wD6G27qAwsCLemiAcYIGZoovcFsUTx7Zh0F1dABSbCzRvJ4k/Lfu29
M5APmVfUOEmUHVsy0SzZNeDiIes05PgIn6o+QLEcs2wi9m7LUmrfWxUXmKK7GR+zSDuFC8vB2T6k
iYQFpSfaiO5uewvM2IY5o2lcMt/oH50mbhT2xed54aPZKhfsjYF9UqVQwBM2/HhL7Zj257AD/nmF
OXeWsCl2wDK7ldMwJQiR94ZyiJqx8qFkYAIROUQrxV6iQo8LhenP+8ZQrDhsQNsoVgK22+yexf/U
jLEeDKOEOaQ4G/8KZvpuktBEcN/o4jlTo+Lql/ry7xiljml/Xf/1I6MJIcbKugGjNHftvwFWpFa8
d6JyMgW2HZzulItZDkJJ/uQgSIsntsLXPIjwSLz3+Utfw2kLIkK6i0+Q9cotE9XiDmA8LBJ3scp/
Uf/YANBK+PCtXlaNF0ppdxjyUkrhGtW59r072lhrRD0k+XXVlprrnwccEM4O7GstS8X1ajM9j/wh
LljqYXaX3oDaeEPuQVP3nXvda8RZnHwgWESU2gWCdHCSNMmiv/tWZsnVFd5D1+o3ma5XdTLHedD4
1CePIg25d9RLK2EDF+9fdWmDxk5Z2i/6C1z1hbkfG6ViIAjOvtKe2fMFgntoq44EA3Z5aCOaNnmB
mlgjO1Os1E4jE8Xh19c3gwKzsrbxMdM2Efj3GMeqTBvcM0Lu/CHlJmI7TTti4ZhCxnhm6IxAZdkx
W7rfqQEzkkqHRxaFlwK0Nz9gef1yl7dWf1QAQUaIunCoMVO+EA8yAf7VCInfn8SO4Wp4SMVAKyiw
hNyN9IoaBcHdO0MUPq0tvZDFn4baVAjpARWmxURekRzRxxhYODQsgQJsiCqDga8dqRJjFsJTyOaP
JSjQfX4lrOIFZj0/Yc4eaIxOmP1+5OyiQJ+8qIhkfZfSn9vCE151fwiaDGP2bMRFZX8OG44gBrId
smFbET9I/drJb460MOAGIfrTKlLt9daAXxHuL3H5m4YxOywqaYbQnLEYma9ELFEZWYuCdYhfl4vE
ePjsGk49Hl2bSE5T8DYANaUXgfc2W7SEqzyljLAzyIauLQU1w0nWYVrut6C0tnHIH/VaQ9b0bZd8
TRmloi1cu+dZKb2PXVuDrNGVOatwWcZpCc0Nf/eQM5psVfDpgk+W+MIUJGwJZpMdf8rWU4UrXAQM
On9FVSZK69pBxIyaUflwXnlAqxBxA1RWmoP6oF3my3495JADywwGZAruBa3nsfINytjKKhFgGwzs
/NysIDC76HSPkfBT1nDbKwrkx/LmuWanhJtWaQixSrl2UkJgY1fhsO5zf6VgIrOe5c4gPzP63rEo
O4RWuH/eoZWG/M1HtuhFxQzDJJAF7SoMxPt2cEQW9L3yh8HPEDJ7+g/x9o2u9bFbPHNn5/64uBFc
SjHmFa0sC4Izcsz3R4bFDWGgn8c/fLWhNIGswG50EMpt1smldDhkwUrQ1G78wEfhiY4gnkJicF0C
L5zhVwQp8f8wQhjTQjof2AQS++ICUDIX9RZT1jGfFF/Dvzi5AGBQq3+hHwsoMKq+KvrFEKm4wNH3
h8hE9LEx/lr4jgLmqLCOX8c3Lp675VUn3DHH+qYBIpV/AcRH82L7cGzb7ZIjG4ST5M/ythkhRV/M
GZJynH5KS3TwdpmKo/eaMiks4rhkxqCmoTuV+uFBx9ZrdTYq4ZWUib6mxEuRqpd2+3aFT4yR9TTJ
V7OJTvb0WzAwjfHSpWObfkEqkk25ULcaTaXDd+EVgAZxp8vRAQ+Ldm+QeTOC8AkHJqMSr0dYKz38
4KqtigKO7q6ncES40sjzmgomMKIu39dByEUMc2W8e9TszwI9au+C3W9R2v2fmIueqCGLd5R0kub6
JLUkmqBaedYG45HfW77rxoHcQCdbUmYAiHbGGI3it400j3eNwg0eIGR8AT/BaAHvQ+iYGJfMm6mL
yWwYGg7NgHOBkaNE2G6Z3JKcbhZToYka9OU42HWLNhYIuQs4en6eV6JaYAo62fgd6QAB5qs1k3ZR
IdhDe2J4h9CjdI2jaYVufWdTDhS4DHlWoma/cDRLIFQ/tFHVw/MfRPPWaVDmbIgc7wWTOTRVri3a
P2edLZ0I5By/QXdQu495ER/AixvNbb5xNALT+R0iatI76unWuNtVZ3eUqQciCrdudwxczToqOeCW
CIpt3pzt1TCoxTzpH1u2py85lY93DW2hvTnvRla2/W6efkqnudB/ln6Js3IBlGciyMWLPsEjEfFv
fykOJeu49B1uR4CKG1k1o8H6BFu/ZpdzYcaRbtZwhNPrK5J+dsOVKzjYcIQadb4y1DYTC6d1zi3r
e41BNEJiBsP0VBmtll3HG8OOgDPzMbgu99xjDhHqn5ECvXZP9rsDQFqLfx4nH39lPzGf8q/CJqI2
bMkkyAgXKTM2yxFszwBrczPCV8XqpsmNF1gKd6Y6lJiLFte/DRkcBvLyoMkVNCvsHKaXDq3ORt4n
bIcdtWuWAWqqqe8lncpp5HF2z4gmQ4eoUDRoFe+JjHOni1rWAVTxMv8AOSlE2bBY1oja9pnS4K0E
q+DBjoI1fgUNnfF/a54/k+YDTc8REzPLs9bd5LPvqrfpcan3a0i2Z0uZJVD75bdS9TBw04R7iyVn
ceSNf4uIhAIqXW4+LIs8Kt8pOOU3gUk4YPDf6bSMTpmjiiuWV/+1mYBzY4qNSSuMjo3I9ZZmy5Gb
hruYB3Ez4QX+6GvIbloN4sY5KASmabNC9jZVQmAoVVBPbKzu3Ab79njaBbVHjPbB4mjqB3v5Ex0L
JekiDdM2wBLaHqzSFh/9QlK2t9yPwKWhMmXFG9riiBxtKrx/erzpn7AcR5NKzsAQVbIoeIoDeyzl
NoY/zo+KTjmQaGcCXfXsIiSImANP3ESJFqu9wHF/MDwXeVNWUgl68NF3N23pdmUekeWmFJVVji7q
aAj1O+VzHR9DTQLpe1YaO0G18AKgZPyr0b6qUxM1lfgfsJIKL1k50SxIernREGA8yddfy2vttZbB
iEnAyPK5sLdZ4Na01ir9kcBntyp3QsT5IAwRZoI/W+2ZkzMdjGQNYnNZLGcSlQQ0iBQn+JjpHqD0
PHUBhPHpwOU4NV9ML4NPEl/PftGx9BOfhAb9r/C7hpvu9w/iMgofEYzwLqnZj4BXWYb5JM/glq8t
foePXFfxy+8W8/cpaEEDBt1Dsv8nfuWUD1Aja6oMcz5acRYn2WleZL2eAxrCt70BDTpRBKvSij0G
hvc84UOQf0WrioAlOvjx5KD9a2kkZxgUIZ1sRXZnZrr11RFlfzVMEQdRsvGMxTtuZ3Jncpqyj8o8
ryrEFUZTsQ4mtwOSG4w9U51HB0cfilrf5nSldONiFgfkk6PvyaCDlcF8tKyij93fcHxbXLf1mzIK
SF0f4wUEsVvkaEEvFT5elfBWOxw51VtacD7518YGfAekyOcfgwWZItfAM6aX8OdQk4xkPrKmXK61
u2mqRAyiGuTC4ld8lSrQl6OER0go31bK+VbaYDF7KA+oidTp8ingKvkV9QX88o7Iv8zuPkPEKJO2
RffxUVj2cRk1it63MqIJuAPOE7HT54iepKNeHJVg2mhdLQDslVnK8T6gbcjnHjk5PHcm+nW72Cbl
6FPFmntTlH/21YlimkbBkuiR3m3/0tYvcVfi2jhwbtB2Hm4D7JRiCFRugJwgEZ0lYhpjZkuQ5RxS
cLFf5mx30skMD1xtUAD/vCrKWZ8E/ZzHT/Y//c8rqrzVxUB9r73IecTsroXxYyZJ1iUBdag2MeZp
M8bdht6bIQ90AQvioOBNj2n6MQphxnk7omobE6d+iWC1Bwb3682kHGWPwFY2PntTC8xqFoTpuBo7
WUY22oxNlsZY2m06+nWZTLDQDfb4rvAzqtnD2mhjMHv1WzUZVyDK+sKsGfAG3zPhV4h+fzKNs4p2
0FdZY3cdKBQP6skQgw7sSDC3TSNrPaB72f/2oOBa+4JGS2YasBvJ9R/ex11fjp+uK5jHdZhnM+J1
DI2KzDoCLVstjCiUD5zm1VwNelDWJwyr+me48XyEVerUo4rBg7Tvj59c5Nnp5+OZvv1EpTGVhFE2
ivCarcA2jvOFD6/+N2NhUitew465yruCKgmILxgIJR8BOgGVNSm3tUft4qc4LEM8MYVOyyCBTlcg
iotsc2ivtCHsbOVOWMo4fwBVvO3ZQVKc4i9jR/TKjVlps/ef/c9f3OMm5ud0M8ebSagTkduqAww+
0NszWxwSw0bbRuSx0PO4H4eZNHDSWGbqGfKx2xxezMOKiYpinm6u3IY3pVqM/FAb7i/H5iUN/9Yt
TXimf65T7pyeXFXcBKY2qtKGMEPIN5rlr5M3xV5ibtzq2g2W2OO3ol0AVCeF9OD21yFP4Ua1FrPS
HrBdQqbpbQic8pIgisIlFWV4tXymEJjToGZPJ6vmOZUq6mSuAwo0Cw5w6g3mrUIqFDv9zaSjFFnL
qNFgKxXPFlSdFFJPolxzAkOoiUdOpIKCrBImyHx24JON3EakZBfjv/K3Y138zxY2XTQx4UMXZvuW
f67xqCrE4kHqt8bOudioXRoAhfScfN82/uvZazp7e3pdMZqLrKci6XJrWi1R5Fb3FqJ0WOnEE3r8
gGblXMVnsQYnyXHV5yHKZozJ6EIRd2ptMcbY6ApUYu1BgUmAektbYR5kCvTNNGEReVlkDn/MIJvK
AEmeTXXGsMyCXV59q+qeSnTKPL17EEwpm0b8oakR7He7qubTmLMOZpXfNcG6hsFwbi0oqS5gu2Ik
dATBTtg7Q2CXrGRZXHNtBtgQ5sddlyETS5Fp3nzWnfSTbFxVb9z0ez0KOuoIlXNO+rYoiNwCI3Pc
saWIpssGbIh2dYzR3haDBsEzryybLWhY5ZPXy6C5AsLoE/otYwqBgJ29MithMJ3DpQmcD2Jv4hEe
gBUKjYfXmKs8ALZ+UoNRqdndNBmzVFZ8ADFeG93s0jV5t2ANa3BPekZyWDhSz0FTC90VlsUlvvEj
a5SBIftj2IIQRbiZe1EbFtMT7HxnU215tr5iBhbGP7ipq7+Czwjc+9cv0KZ2u0ZKjGkx3EB/lmvd
9lHiZLavuXfgHifZ/aOx7UYxwr9xAgPdKhXmFwUfaEQTKSbqSpXXYltY5aaM5k3T3naiQlpPsXMG
0ejZeR1N2xoIq7Y3uTNbgKkNEMGF7OanVjar48cTSRxn3oj7nlDSIIjUi3qo4VydmoKDwVuOT4w2
+xYr3vQCEONe0fReQcu+9R+VnxjEXz3GJq48gMPEw0ulRMkzKAAZxFolmQHweBwKpFQRpAhmFjfW
qwSH+4j1U9ja0aa9BjWbdTe/I8nXrz4NV8WmdGMHznIlYwVa0WvbJjKZf0smTZmKXLoXEQeabxEV
KG+GyxSyytL6Dd/25/7Zox/RJVZhIOqDRwOgtScHR/dCN8IIO5DB64ocwFF1Ae31a+scZdAs7eyR
DICrG6+yiPuLABsXILk1ieIuOZ2dl0SgwZqBB15NtNQRFZ36eABU45x20aCwj2JlDo2UuJzmax4a
EXnfOhpZLdN7mXdkEzBxwI4ukkIekIzA9doX92g6khpTT9rVjlW4qpZlLIwJy1A261oxveZsZIsO
sDz7eKkem3RvWYNJX10g19lsmOgmZbB5z9NZijNLWWyNzE+/B4wOIC4pNNXRERnQtBZFQFmTXhz7
76ZL/mmUccXbVijntb3SOLDR5UJLQlKy4TJkVwJl2MpWKsqLhwXVDwc6N49ik/I6J0/jZcytgW5f
T3cwgeGiiCZZIJew7pq5jMFH4aIW0HpPoH7y4hz+4fWFWpnkrzQ4E1mKe4RFyxeq5Ms276WJdiPt
x9UIoKbn6EFhOi4O+OPZptfHtw9HKiLwYkZDzDyWMN9+7oXxbs2rUaiW3p4H4I0uKsMFnjQQ5HZM
ieu/8V/RbTclinLfEDYFuSQZF3jVaF4iGO1TzePeQvUgBp16PKAJCMDxzl+ERVzoysyIrJwqK3ik
U9J7ZHiiBra/D77EbJuJXjqaP0XmdYcknVN3oIdBOqpiOjHuBaYYWJir3sZzeTbT1ONv2ECM5oon
eXOi2zsfH96v8deUj1XhpnhxQlgn0uo97QIye8irfz3WbALitLZ8KHAj5j2FKcWa7V5B1shtgoiy
SZajhpBqtiA5JGrw7M7DRKaP7mVB0zcZzuiHhBg5UcPdW9kwAxvPMga5wJADVk4wXUQq26TzhPhc
G4OITpgzIetfVNMncIV4QC65/fh80I7nK6sCn60xEJih3eBMLNO/4hPtO6TlgbiBE8h9zhbppjMb
z5v+0vxlLsc+xTRD0TqiPC7LQ4ky685utLNMEyBOuh1Nz9Vtn5JckK9GhnvmNZqu7NL98LVfqspU
vGNxFbN2uQnVE6KugiugqnlnLY/VbOOTeKE2tZ/OmHIkifLHGyjwyePUqAAZHjdkMXcBZHyiCZmu
jtxclCH2HhPNV/V0RdaPhdIsqxawoHNlvxvwyaynz7Xn1tdBdfAAqnxSDQku4mhNfJ18pgqAbFuP
A+py8zrMdTodxULIBXlm1f0W7PzRSPs8KZKaVjeaj6f6UbhEL3gjXokbxafAE6WlIuDsUewM6DPW
NhtPH35220Er7UNqux6SWwy+yGJyqiFWLsCNNScS9VgOeyXLuPJ1baECr9zK50kahRc7ZiSgQzWk
+Irl2eXjg8Xdru919h3xOzTl+4oCUZX5x4dWPBqlS5SnTi2Pm+qpZSXcv6gLbWhp8RWX++eqgB9R
42a2dPNqovf9fseZ+wB75XvSeddkrBSuDHmbLOn8ySCfNjN7D2q0LKhviJmHCEOyIkKKi8r2oEdg
YYL7h/lQrS4vy/u+HqtLkArkQgdId2bxIde/F3p8ce0YW803ieWIxQu/tOe/teBColRMsnPKnBdv
Ghm7M52Hs6Y/H32qT07lWhLjerbVKHujMb6mBKB4bDEhrNBiKkj9irEBYH9rySJR1qmMZDnR2g56
zLaPR3YpRpGqFE1ugQjzWmURb9PaA3PC7M9tIzHcWnSQC7nP1UG7frCH1CZHAwfCKQNKove1Dgsy
587Thu+WakseQ7PboYmctNHDLJE2DYvhF0ZuR0lgMvPsTxVKT5my5/M4Lbc06vdh2XdyXF4eY0RF
uj638r0FqjtdpFVHlzb52f5rT6wJxT8nGwxdRKtkjiN1ppx02g1WgLr6yF60WwowwGnvVpiCoSTH
jtn2JWbE69b7gVuhEXmZoqJJaYpMuORO2p25054cpAUivfSoacKci+OM9WhB3AGJA5IJnEd5PdGv
XmPN/qTP8Z7Ljl7OX45XV8842GHUaABBzmvCyWq1xGEokzY8a95BSw4hJv5qo0ec1EltmD7zmKYO
/C+Y/5JZ+7IAii7y7uAcOPbmKuiG1h/23EuIGps0SfPjjBg5As6rH+cCqNbA68Ux+uTJZGv7gWuQ
2UL7QzKqLUojerZmliH7fJTKMoxfAYEGF9Z2JriMACjAm7wUC9fPneYw/DHSxAIsoG8segdzOUJG
+ryA90VIytWx/yqJGBdUdP6ETGiwOksUUgbQ0hsbJ0LywwoTadNSd3WJw3vTz4HR7OeXcUctAQO2
664dIb8EOq3ynuvwCa2VcQjbGphG+9DEHuVdjJ72OmSjIpt4h2sBFenLE6pO92VchRy78x4nSdz4
0B4z2wfJt2jl0mE0306erXgjS/oBJ5EKpSu7u+GC9+BNP4QexS4fk+3BVAhlyLTNJ4Kh2bzpX0Ez
FpfqnO056mU7tP2hWnqy55vf6xO7AU/T3NCximqV13pey8k40eGSxC3NsM2dGtclZYOc7Jc6p51b
BgcdOxkZzGSppj5RJfJiCz51efw6CyAn7ySYLvNl/iFIUe/ObLldU97hRQ5Wh5Eh4OveJVW+Pnfi
MmzXla8RiER9zz1aWYCxXK/4syOrfGDZTB/YefdYQxI2fniXtMIRbjpAAwXPivrlSwq+JMjv7NGC
Lb7q4TVe0XYClMRL03kKzM43elvHBZL86iHIPmb5m1XGJiSlM/XKSkJWx/mjYUu2mkOVCWF7SbI+
eKCoXnw24utcB23ihBlzDsrudI6AWsNylE49y+6Npyk8+faN9Xj/VpzQcl9GNI10PB7JABJc51eb
2239qffwU1PUbdYTghpITCGuLbF13ay/c/LwzgKSXPVbOg072Lwo9BT3g5c+GvkeeTb1G0W81fjr
pLZ52HPZxnWKQ7xwqeDnAl//XCly2MIjr6rQ8FB1XX0buBnZKM4rvQK6NDCqNQDkgdCc0veO8Iab
XLmGraV2cTWOFUHFAQN6oXSMPlLTUCukym0wneuPUXRKyt2UPWRNLWvUyUHfsBWG2gpD99JUy4RH
n6RnHTR+sIJSu6JHlCgZmfx5S3XrDsqI44O6LyfNhP3EXwbVKsC5bd4jlQ3l+XVM5LaHNkVi3HVL
tzqrHqP8ULz232PJSYxQwIyz5Z5cx2Iw9GXBB0WfEtUOQcWUPnyq4nKVdNHHFKtjfz3BPBp26qkG
ZHuR2hSs5Xg7TOiELtGNkqIDLk+xZ4TxIDgIQNdGYUgKOISRpWzuhpITc0xm6CZft36FNrENg2k3
s61kN038YhxgbSeEov+cAFj1qNUSDa8LybhuL203q7zvtcRZQH7hvOcSz65lp/H4N1Hnhpg8qpj2
+9sZ47/b43IbIB4jtanm0rn0rkVUQHdMMQCD5+Eg1C9kAmXmHgOsfsyg6rozS7qJ5/xLo0damzhL
j9GeS2P2LOdGPMO5iUylWxYDMXLG8xe+QdefiQ763aSHU17oiExAgb7/NmDimX4BgzMXTbRhno2N
H6FjhEuIB/bjXkTy1umGOxD1PN/PgvO+RFl5QNIdi8ghKWzT3RCcmI8JhPBP7WMba7qfA8R3JeOA
Ja0kYL0hIqXKzeJf9BX9zMETiSBsAyu7I6UKOAlpdS226CO0mAyDWPxX0e2JoDmyvgDX+FfmfR/2
FS1ss+9C+lwk22CkOuhUfONdtA6FZmot0XpEpLx5rDesEd77IZMCwJCVQ/M5zlnbgUieQoCTHQ9m
nUW6wNWJroLiC7qTsh342M0L46Yy8DBJlGtHxjWuvre7dE8a2qgXzhTkjPk8TD89jWqWbUiyuyuh
EjiFc7el3gZd0ewMMziEh0k/dhC+anbsryyBki4ybO57v0qRHEFueEgyKnHIcqv2KbD8T1bntfhh
Atpr06HIWfI95ENPtJBT8gu/alomzm+1EaUILmPtwWidXnGoyYVq3LxYNK9WgxuueBwiib2tXmb5
lXu6+A0Y1FPWeNjEfaoXUUyMjFbX+nTZz7EfscRF6JfB+h23eNCs7bTikvLytWlfDJvN2rNEAloI
Cg0ugoQX7TRiHEAIXmC9HjuxEL+gQPCiJmz+MDsh25EVOVFoKvF+CpamaU/29E/f4ZytUkJbadcb
9h0UgapVl7e+YJBxCpMZhZW4Mb11J7oNCCIsXx7CX2GKFJv6JUy8/49jNJYYDebFyZ5yWa8SLwPa
Vf3yxJ0YzK+arLo38bYYYzC6lMsJMALLIZBb5xdsGb3W7dkrMWuhNOEvV8Jq1suS/K79U8ZltwOt
DTH5XoIcJxvR0z3Ih8fi385ZkG40dI6hlaM42fgC4pPq/hq9oJyIwK/wHYZsfyMDepq7ZMfahbxM
w7yziAHw9ANKmqMUHZp71Xa4hmZVd1CdSt8QpSFedKcxMnLfYuoPsBfLcrSSgIOIS6so1DCT+kbz
aVBFAjNxd/QAdKQLtgRyUKsaP+AyfsmQ0Ko++FeRNkNrqN/ThCR4EFKSeXN7nyjeHbqN0Yl5MwEH
3Z7I2pkMdSL9kACD5S16hdZkh42OeOLO9L2KU8Fngw31EbwN66fLj97tHLnEDZyphpNzBBkHGf74
wd37vWYXOCtJW0+kn2He0L7ARYOqTjG+DylNTNjB3CdJJUoLc1zX2hKCL8+EarNyy2q9QME7H/X/
FLHhZkZi63sFnbmkpFa9AXjcMNBnAP3KkgnJXkyyoxoipO/L89LTLDMpwz3uNr53SaxVt2JfUPl2
viFV3PmMWjVNf6JaXaGMjKZ61XoUlL03BQqjCC4elKKG7bCc9r0A+VMe5wUYme9cU+9umu4zNlpA
ORYZRW1voM+THo4O9YxU97n+gQEv6rU5Y6v8JZrZ7N9hIDd057C2V9C4a3HyOeJ6OdJ5CAzdl+yS
iGnLyTfzXf1drKYQAdagVYASLPmgJGGk42pkBmUnER0h7M0Ss5Yhr69yn4lvQCAHsllyGpuKvB9r
QtLu5I9IwgQsnmN08QUT3MFc7j7Vecles57K1GlYs6G9PDqjWqou2SNQXynphFwwHKk9rSESVTqh
QUyC4sAhthksZ4M7S2axe8qXWzNZkG37Ggi63x1OjsvZ33qfMwEu+p4hLMMt45QQklo8dHx1ts+N
xpQ6A2JqiV1FgyVktcGPoLwVQi0B1Apv71umrnHJrcUixQHp/1uyzuKyljB2JMETazM9V+MOpDcH
LBhwfNnTUUeXJXbzsAPk6wSsN8YbRZgIeDEmFYhZbgi4sKg3WMU32oTtHsMvGh+ndPvU70Q3tUj2
ZQvoUuS6MDcUZIj/eh9AV0y2YqxZ3C5iY5QROdX42tC2YSs23ebvsRw6D1ha6rpe9Ua/1cyQWTgx
jkamC9uQZ/h9K0cp5jybOVYoqvVA0pNvk+806A/vsn2QT6xSbBrRDjdC0U/NPxKxWoOCGUk7sV+B
ZygbT67pVgzwqPksHJ2R+BtTgAl/X2/knV/ZA8giDWF7m5/lvmcZkKuYV0Dv1jBqD2SxFz9+70ML
YGVIpO5gqAnWTJK+wY4UqJs7BnjqSrMXugBSQaXZYwp0p2B/uUTz04kW5X6x/eBQORIZisgn4wLu
IZVFI/w21qO4zP7DpPbsg229CfO5C3VCpT8EfKReIwgIDiyLdo2LrqQFXXNSG0JgWNcQ+QYICwL2
SV1hrEUoB05veVMDxgEbqM2OLSNnTRwcZ5IqsAhy+NRL+8tOkrvMwonbVQI3HkgerW5m81bVBceb
+0S1oYeHT/wBR9OU9EebXnRZGac8O5aiOmtXRQU68s4LRWEdxZ4Fe9kumcEKXWyVQoK/U/sGjpsX
asF4hKJex3+5tNBvBkOb5Z4IAc4oIRjRaSdT5PdOMOqip7YlFWdaLpcuUV0AdcxjKhoN2LKpfKFt
YHlfPg3bxDnNr+Kcz9kycYjp05ZosZUPq/95sZs28VuRKUFfEaPWpWpWGdrHj/BzarAntYaJLBHD
qcfw0iJtarPf9+8k3zhghlEOduMHaqCEIuViny+W9OLVv+37kBszAtCXX3bHdMtrxnnBi9TejR9G
SYdpZlpUqu8uA9p6Lqf9ZlW0SIFjYnC8aoXDjCMVlYLXOkAUzT8CHqeHbgkYJapZXDA20iJJMxFJ
rIHw5ruPqdLO1GTe7eCdEomAF3A/2TYpvedWFAH6pFkawlumKh25TX6rPDa0Y5/KsIVFmm/Dlrt3
lykbTO+3FZndKs/89+88vnnObqvi5H2/LesB8PQcBpIRBKqueH9nn2othjyKKFcTly4DoUVCKJT0
F4bdk6C/PZskMTCIWt/DaL9zLpvcJ0zSNTXro6zMGnztQQvtYik685NcUpllrLxpu7Y4tIlG8eJ6
xNl/NNXb9jrxgBUCgnA0UcgwqpoLZ9gcOgRl0Q+W0FBMNdIb0sSF2rDvbHEeaIU7TDj6lgmvMP7l
zV3JQRxPqBC9fbaNR0sqhTTm4+lkUWNqEoj7AdICAlggF9/nx4xYkHHRPPC/XL7KXNxHXteU+1o6
jmcqwt/GlTUe0Nu1eLOXXFnn4MxrEuj1xvkd5yI+eDqsweCPJXfP4g1vkJ9uDHD/GJWJbgbfbKqn
QoeWugm5wOSjNQQBexxBKaYGm3Ed4JtFYyXPkPPXkiLj2mfjNSM06ceKmuxolzFld6FoQPpa9eEw
fJwMqoS4A420gcCxW4tulu+HNEAuLPSk0aPY7kHgoqv3/DYQ1jHb4qDRqKk2hb0zPDwyKKr0sSXM
YX5QeIvkffgHBKqJ3EjxgMof5KvxrwLQaTCB08jZHUUAxEVvVX0G/l3C6bCCrqYLPLVijePURMtn
cPL8xCYxggqD4l0bbVr19IdRFWY8ILtfszNaPRLMuZZvY0KWI/tCOonr40rZwk7FwmidVGHrMFN2
Z/c4W+MS8/4wXtKw8tMVQuwCV7rlx5LnllKKXIQjtUPQwxxQoreBRABVljATA+BSeVT5A0cQoMl4
CZ/y+Wv2J4TnFsTLe8JjPxeb2yoUta5/InmT4SAn0/eX++V3c22PwZHFMPtY4yE35dGKmE3IZnbc
rUwnd1ueboxWql1TZG6QmIYMvX1E4P4tsW+ouARjliQQFJJP8V+wNF7/6oG4qoN7WQF6f7YTMAn5
BsviRD1mP6USFrlDfoHUK/hBWpxVzVKVkIgBLBiQIOn9YvOX5JtOJ1bzxrk0MkzeLkZ4Dgi2Yzjj
Fg7qx9W9TmoHGKdISn9TnN5/31vkCYxMhTXFpfdD8PMwlhm4kAMAuWb7KATtE1N1Bp1tA2EpVziK
o4HH2pvWxKD4UzyYugU3tHAe5MP5qSjNrPqxyGcFs1Ah73F4dA+VizaBNGp524izqo9P44c3Xg5L
SYmAiZkuuwWErLDsFdyBBUxNJh2r7xM6PGU4h73bJtgKrNhD0Ylixp0MB+wepi50q1VWm7Bcxfpn
oY3Wv3xJAj8ehyf02kZa4i1GxQmzJ2p4l+gN1bZbWtCOFGW92fijehlt2VK/jhg9kDMFgD9hdtk4
+NWX8zP6abmHo6k/TZMZTD9NG8g/XwEq+h6Bp2xFTiCxtLddogxSlLrLQH/3fWHU9g77zBB3Z2ng
fmEHs9ZAT+FXgt0wlTtuadctFbLOLhh0GDtDn0JkfJ9DYrc0EvPI8jpNw/RKW0qtyJlwoZMjGzbC
z3qhJDR4bRp+OvMMicrFI9A9oKtE/fNPQ3LK/70kBpZ27UEh32M02Y2p24OqRnYhkY2dycyukyrp
cSzyu62xqDJXVclSEEmaDbNB9mku7ngzuCFKkX88OCKBYr1ZkmAUYTmq+jyeIsiOJGIpbxHddqUv
p3lFUpWhzLDVBF7rsybsGDuFYFI9DYYf/nuHnHRz6vUkN1g4rrXnw7lHNWkD974m11wybWofuD9O
KHCU2jOU9wCVzMo5ZV2u4Rj0J0SS07C6EzSkGmY/25J79eJ9lE/bFlPQjjbqOguaweTcIg+Uaavf
igsuiUnjb8AdCyqLZ86WAKXXZqq2O0sPQuTRPBTsiF7VMPan3KSEpF2FUh0R14O5jPyenyO0ac2F
ns+9mxF/kxNnpRJL/AEUBJzM1I6+0tvZvRXedPNQt8eXiaIdQzGIQcrhZzT3CnilWDba4tGdvTNn
XkPOInhXjk8h2FuQC6SLi6UQ11uHmowLTe8wzwfCUzNNG/oEM67MfjKJ3zfxn4KcofKSm6Rb3f+i
DnpXsjm+bKTkBZWEGyfwrbDtoaImjjnvjJxvykOWLAQVHrH1AQluZqWTr4kNea2Tm/f9cVyAxSTq
jZ0ZBQ76RhORZlZsby3RGOtvkGLFXnNzIDrB4YZBQEQL5Gsuxc7yPbawl+lQa/fqLGIP14uh9mQF
lOS6Cf7cSMz/1WxwkAeTi2Y0M8+MZR/Lz++nPWpaOkDB+KJ9WIE7fQ/s/D9Kwh3yORAr7Ouba7Sv
mKZl0TR+DCdqG3Ogod4KNqXY6w5Z+gJB42i50kElHat3PcS8sPZF1rdkK74UrV3RwOQ5xXDw5qxk
UH123RcTOhSgUmey1RX/BdzwpchaGpUFrgsmt7JyaomJMl5zKphBdijh/Sn5yT0zZhSYFKCj0v/v
Xlb5FvsJ6ZQwgMGwq4TlEyGzzfZAYAG2gM+qEvLQk9nnmO/iPWlRWXI0JzpbyUQ7aobz+3YrqiWO
vgA7JssKlb9mxODG8v1rhrpHZGP2x4fW3WnYneS8wVFPacsyKkaJOFvHtY4eYWLKEP4IXUl7Cmxx
pfgTFasZR6uBovqF89b/t5FR+94yI8JX5HN/edSlxS4tE2QQdrsS2lXuUxdzra+tWRo5LzUF46CJ
LxDbfJ9r2aScIDRS0T+O1SpSJ7z1v0JRGJ2tu2LFTxcjLfEp8sxAqDJCwRi7CnB4rkfdKyt+A4ix
69Q5XaYDY1af4xfY/ME0O9xZG6DZgFIR7nYE42aPHhbqxDiPfY+qAei8NoMCv1PRn7EVZDC75YlY
uEVimEMR4FOptIIo6vZXPhQvdg9X89DQvMoqi9vSFwZzJA4HNg06B+EXU/+cHGPhsX/Dvce10aDZ
th1cKVzfK3F5YnfGwYj2NOpG54QaSKRYb9+EaTPe1CESf35EzShQymeDoWCew1S6m2cnyQX4YGF/
dbvZXR39Kxul7tDFpsAaDoZg2lsAebTynJXbEvP/SlUyiPMfE5GG/R8dsyKIPngl84g0wMMVAZ55
7M1+c5dAmTVLTBPUUNOJE3w2bpuaJPu28ZgPigPtx78a9tT4mvtV4kFLGfd+0qN1ytzyn8ijLAp6
SWxGD9BUyK9NSIUOnXh2auBxp2K+I4Zv8GJToKDuPftcB8nwsE3CdNEXRo6yALZYjHG7s3cQZhLh
E4IbGYrsz0xeOnByqcUBQxw5XqO+u/0VkAkqRDY9LOu105bKi1BEGRRbz8nhSjWbPFVRZPnthRmn
UgUxmSip1dTpdm/5z5deWLiL6xML84tMG671lW4jujFiyo5QKHhZc+6Ix4WCjpivXv8IpPm41ADu
eAcY18PJhzY5+Bh4fkw/lk9RujB1/r+gkGhSR1TpTcxVbdmjewF59lG3kSZy5+UrnQqo0WxUnIPi
36PB0irs5FrwPpw7OuqQtj2wlaWSUXSJ8H2MyHNZ06Y0qOCczmhIBfiiKLsvIcx6lsbQRHWcX4T7
tInRX5u7Odrc3Qj2Bmj+FeK1cRqS3YgTzuYaVlCpZ9JBPCDQxCTzbcxQ0tsZ5j0b0wyRr1Wsalhq
8lt8/o2e6w7AmuyrsKG4nXm+elfiTSlASkc6zf7GUSiqRJ08Wi42u67kmhJ2TXwroQxcXF+L3qkA
VE5kYddrVSBKVcvup3gz+icvzOxvpLTg29r4toYrmaZSbB9h2RAGN9+6DhOHYuf0P1JWPCcxqk7+
cqPbQriSY6VbYjoZdv4FHt1XkN/ivhWReMI/StjtYz9vEjnhD+W1QOUUF8FkbR/tFKqPzBQ6H+L+
WmXZTe6ubqNX+WfQviASv8oJY5UJURhEGutvHGhUuOaTNjUBPYs3kOaPpI+BlTUToHUUGcgxQ6ez
tZnq726fjwBYUqOPVSBvpx6iyxTLRDT1x9JAwlNIA++aC3PrdnZpMNE2H4usdBtvuvB2FIi4kJ6W
ueju3AHeTCfBfp8FSpZ04TU6rUEyEUjqTVJQxD1NKre9PfqglU6f4M+ni4JVqNZx5h8SzSiK93e+
M7Dx9fD3eyMKItayTMBkcTH3gQ4PnwBIVYXbyA7ydalTDjiO/blHlVvrWoqIBxkswhmy3fsXEOKl
mm9NKKShJ9OpZafu/BnvvEqz+0E4ijS4XOXaaTA7BJVJsyH6Q7/3O/XupJn/2T5KkAVnv2b5i6A4
jh0D/PWLTDrWKfBXHVY8YZRsWWRp7osQuoRLmzi8zexZEY1Yhauib4DfdrjvrZBs4iCkSxfAsjL7
IMLuXLKGKd5M1JJNueaRjaUfiqCg2rUY4EnA+G8upgWbBwegd3zjk9em3V5tHoa5FDySC8lQ/cCs
nwxA2Gn50phPdrDMyM/Rfl+ntzSxlRl1B6LwfgPFz78INFAxwfqkSSp+xaqGQ8Pgcup39UCMU74m
diUhopLoV7A91mnuRnrCA6vQRpOZju2bDEQudC0Xri0DPdoawpNBQ+idMbf18IyHH0v70Iq0JD9/
hv5Cnr6ciB5zdhoPiB75L20s8CMmYx97bDJJI+lfy1icnYQuzEFHgdl96dzm/wfHHDV5Yfv6iJEd
a1wgWWYuWCLxAo5FtTR0Vy8SyG0V4BR9P7s5ThQnK4KdX/hBYqN/tyGj3jcp3a5lE+vI2qWs0yRn
D7ihg7JvBmxAATJqWkt4Ux7OgVrQOohZ1fJMjHKeK+d1nDXyM7Jj63Hvh8JlshkmrC0503qB+T98
g3LX3PrVPkZly3CKtkmdobi02MvUTbi7IIdfer3zmMSLs+wsTcjdpC1rXVdli3n9D5qECuwUg1Rp
/ZbgMfLwuwIFKOl8a2qD77hcIkNpyxD40OmQMOJZjlhe/AMUR4fQ4XUI+6nyfoAH9SQVXrmVE63v
KcozoO8jwhc0Sw+4u3TJ9nUiPDRUTbN9VEa/G+0PSVmSgeIkMS1xFYPCMxs/j2JHA6kMg04248H5
9ACQC+C5vGcGJEC/aFR86gW0eoY1HvYjHsIG2eSsB3Tt5TbjrUb7KhwX0e9ROP1p0iv8pWwA1Vdo
WvjIt/Ogu6C8L+NcsQGbMpVgww5PamObd2444N+Lhu/V9Qv9gj8OLvhFWIkwdcwAo0Izsqvxd9GE
DK/7FdAn+K6czNq2JfGqU06lYVhGS42Hs0kdD9jrdBsU6d8iCQPZ5jlDvN1GwzhqL9COChicsxd3
2BCjbTK2I3pndWDm+JxUU/v4OUH/5gpOBUAt4VWEEtyayy/qKpRH8QdBjazEmDh0SxnjBjddBHKS
WDriXzzROUdDkDNABM9aJaOMRgf4zSIjBpJJZ9be47AbzcY688KBxBPeAC45SpYDBBVoDsPFLv5j
hpAqPtRwzVngr5ByppUfrlwPtLwzeN6X2AjJ8NXX+QnoZDi9Mcuyrfrd9ac6qrHmXXMowOjzSm9G
JmiENxgD8cOGtDnLuIXS4Q64OIjNMxPdQobd5NITRg6kBMEkDxUsKZ51lhnHuAgH+mJp1kkSkKfn
X5AqjWktVO6Gf9zHXfY+TyjcQoGF9a1PxP0jE/XFnIw8xOF/yxZOYyKmhgyA/PoiXC6Xvm3b4sW6
P/kOv7SKzv49jqSS5r/D58R+AHyOzo8bppgL7JjmGscPsmtgdx9CR2rnpfSQOLj4f+7U29nc4Pq9
eN4fHXZxqx66/aDI8o0RxYNUJcqhcDY6hYJ2yBYq0baeh5Z8KV6eXzQkcv3t+CR6WmABi30D98RV
t6scpu0XqkFqdNf1uOlIPDAwXvAE/2HbK4H7GlToV/BwwSpZJ/t5zKMwHgkSyHiKCgd6V/suuNe3
iQ/sQPgCrJ/HCQkiF3Xh/En+N7wKMtjJOvtnqFxB9JtRoktEuPB+MVwSQdEf3WOb+JAJWldl5bNO
dDt2IKQxCICzT/MwWLCd96NSu07xcGze7KG+FP3jJeQM1IsT8SW24TEFTRsVdCyxY3UFs03YioXy
lCgp8hlK3MfP96z8Rk5GypcHpttOTo/sO/cjoT3vLDsEaNWp2Znkn6Hx44lHsYTcdnbHtNe7OOuq
KSqETpI3iS1YC75Gm6u/wM/MauSpSf61hB6vkguMsOAl5VJvnrg/anWw6ONeH9QGwbwNNW6/S1gf
Ar2KC1yqdBncraJcLUbRX9b0giSFLxnjcO8rJrdfoakgGIIHBfqIgKfPKWVRgSfxqagquYMNck4W
fK+XN3oQrXOPbcVoiZBkJVkW9BZcbdNIk9THxZ13atwpY9QIoGfguTJdrRww6ALG3mSWIFRUXZ0J
yhFkSeKzvw0h0mSWh3R+ENydjCOCS3IqCwGFY7fByL7IUTMQVSTkZw50Ld2T6jEU+wm+lkhSYc4y
/33LTgAzwIDGpgrEcNif956M3/Gx4RBwBvvcWB+hwKsbjW078O8mMx54ofh1f3mtHUkKliVfjB/D
voCAzWa6Q+Fc0XIB12/r+6qDLLfN92hBN5lI8V5TKKWxYZUeZ/sjOHGP7el/iwYSs8h1tpARzLmC
yk8eVr3pHV2VeUpGDYutBvYyHjDHzsSFIuVg6/uHpVZkSDPqaHovaz58xLExCy/6qWgpLYfEBkft
uGZk6e9xQG9chIzpdneXD6qH2x9LCucmzMDZ7IL57yUZ4xhpXmX6bEOVEJiXyTE8rVbFj4+orltB
I7aTM1zIxJqcmTcMSkj4UiLy3zpu/aABQ+2jKsWIkueh1qobzy+dW4EyXZaRpMDlkWCetkGM7Rd0
UqynAUbqgA4O2ffyztpLXmp3bNYoshhp2dOSBSh2sBFE2nSUnd/zuGdonAZYSlIWMaAtZLpljjmU
JfqdPPDypAbfL3MQTrMJBThHX1XbcXBWX2/0bLtn2vkVb5e2agV5IbUP1dkIavKPR/RGudA3q71X
RmZbRoJmhWxj9X4hhp7LYWB5nqU+ace/z/BXXz7d0B2KS6uILawf0/mP66UOmhDOPTLDd6ZOFgF4
29xtdtVcPmOPWduoG6zAbZ1h5pcqop6QvmUXnW0xtklaLU7p0z9GNyStOy/9zQFxR/YEmXFGb5LE
CTaAwlXGbfOJ6ABXvfdzu3KJAWpsr2xkkT0zQhaeHnzZhsaLSxiTMMbzmzdxI6UuqUsiPbinD/8j
m5+BbGvzrj9b7YJU2ureGynALsxTnvxf3FFTKknP194eTPraoWfNxaa3/V+Dud0HumU8gDtfnxX5
leKFmenQRIeUf9oA+mXQvwyhegIVL+cdZkSR1LOGiSV9YztELuig6XU1ZhbL1m2YIeYqYT54FfGK
p/RxofCfu5rhKo8jquefljwgllVxFvbj83NPP1iEOnc4ZQZEFlzdYPeVYxwr+c5ORg3ynZdh4LQ5
HO7Y1kVhYRpyBQMYlghCsnJOb0kiP2oaAREOT5Yz/Jf80Jr/ybUHuzqWkM64EsEPbwwdw6kc0KB8
D5oKgUohRUfr4o55S+9UG92Sorcwypcbu7D2x7QI57VGtwKW0zdpT3+AtqLfDfOcjHe6vxkZx7ja
xDAzf0ZXPYiY0MzrNHtwRrJaorWVXNBWpdZYfHk1YKIZh15dBk++uTgdR7zWGMynEnqan8KmIp0G
CKYRcQ7eKrvO1kWPSfxcLlCXCOENJt51xSIRKgU/Me5nBml7NLJDJdLhj5NE/R3xnjuEaYgJ6w1y
Pykboa0Mi0RFegilHD1KVBwFvprprzaUbK+Of0sgdbizrB9HqK7s97RBTkyy4HWBwNTnydPtCkF4
VfXFnueKXHRQTvSwpYqifPpJzWSHJH0ALaRfdoPSRn0e2KLdHvnxY726MqqlR8uEx2bimPjlg9dP
uIT/F6y4FqmZjzFO2eQSpEfJxA7CXbrkleeOfMkru0GQ9MgrkDeUrGrO2uBXMHWtqL12jOpWcnC0
9NKzC9bZm/eMCIvf/gx62A84ZU7mFGGS9w6WTUbRjH/B4g8AE5fHqOxKW3x7DpYYeggOkyvPfef4
2sf5Ka2gYopvj671CxoASRCB4vSg5QKEdoqxdoKZfPfL92apIurJh+8bV07C7KqS7fDDSR0o1XZ3
QC1VVBl2HUa3bEtzuligwCmUjDRmdrMYw2YKCmc1vpOzL1+w+ey8e/XZKIZT1LPY43PfXFNJImku
WlTr+niI0RkC0RT81A8Po9aowUBDVdcM89yByHehnh4sEmvhuq/prdGAjYB14NlU01mP76Gjq/in
O9dmucwH6vtd8j7a5uQQ7d8f2YICicF4LiNszcS/JPbUyyC0mu5LFvOlkqPcj8QIWSZbPzyJnUlt
1GnjOnmFnWj4QWMgtBk8ot/9nRpoGdpcMUJCUkPWzokkyY2zjY8Kx3BrNiMby47lPJKm9FqdDl23
Cf6T5IwedCPXBE/Dl0b4qm6R9et1H4eNacy3fU6z0Lwh28YxYVorZhQrqOqHSBYZlaEHGnMxXLGx
IBP6LBAluRqjmCSrVyMxlbq/j8i4zXGUUIA2R3picKpF5VKzW1pqMVWwsIzgwqxz9M9WYvHKnsAE
TiobmAxpMobY/PNDZU+uyehAxRV5lLPfVZv1MaRMazNVN38GOPcLbkjgEn/WGkmYA+LbJbM7VS+X
M5Af2qwirmvrYd65Fx1pgPK7DKWBJxIhpudG+NzD3uM3Q1QJMeTMGyOWXzpEkZUmZzXcyOinl24u
CtUiPcNHu2Lqyc3J0WvoDuwdWvxredtDjatuC8tjwYlgjIwY7FqNRpcir65gCO1WzORlUKAPQE4W
+ZgzHVTdtzwtUfluffnAczbU7zTuH4AQqMRvhvJL8MdnLRtPHGIRvuuKtOjt8XLgNOXfQsHpZYAK
7ogIb6h0AibZTJPNxlxHQV7n40Gs349uvmInDKbgr+QhqXFJdbkVydNZESFfZuK5KZrhLWZ3kWqg
LsNLGUeswHXgxYlAnxNNEYE83NT+QmYyuXTkN0A+zlN8hDtL9WW+P6dH8F7we3fELSiudyzwcgpv
gjIJ+j13siGMOTKlnWlzVCt2hQj6HNWeNBD+qNf3pRukzzXlm4TdDQ7yVrpx3iLzO7HiWqHJdM0h
RVpLdVO+pYQN/uthXN11B+w4UUO+G6udtUzXGUGf0DAaGT81qVTwNbE1jjsMJmgTLo9bX5b4b1ob
c2/TeH5Z1zUp2hAiSpkv9OJnmBHjeI4NGalpeLygRWoWn5x/4Y8zDAthZOhWk/mNFGvV9hZ84HNH
vzWogp8TwX5Z9mkhRBYtdPIH9976S/+XudV5whVTJclZVzUz6u9Y8mEmz39E7kXM2HzzrMfUl/5N
notNgb7oCmyKLckZeO7J5Ec9AOOofgDDDROwOSx8IOO94UEkezc/YJtAT6/e3vQL1vbosdqzmuKt
Nq9C68Tzd7vcYtrsbjG1MjUSIZX2DLsh6TgCBgvcrXlyzQ+32uXfRZblqvD7ftQ1hs03uvT5U0f7
HvsZFxifP0wTCL60jMvmo1R9IxV2Uev/CX0C95MtbIGaoTRWLzvEUpNxSIkPXZWVrrnDzSQ0uN68
u0jCqY49qrlav6PhaobR9AtssNjHEfdg66GwKJKVWGKyxR5vOWXvdcLTW3lKI0v6+MnZUR+URmzB
PUQb2hXQboSWmKNNts82ttGpVQvZd+tx/bQWvy0B63ICfRabTBb6QsNjU37UwoCLwnvHdKU6hk6n
pj5gzhouQOwRHeXt2xwQRuvJB5uAyewl9cNTRMsZICPVx4qhiKMA0u5vyydYxGmzCE3Lu3Scl8WT
yM91pd8+LHIria/Jn76gNMbuTeGdXjTV32BKsVSg1hFAqGxXYPvpervmseKxfZCT7s5mPlmc/wcq
tWnr2lf7KrNrmweosFpV8z2jYFB46i9GBd/zHaLNRT4XR+Aeguaz4bnmKhpt2Mg5hhWzixLkkUm0
xQCRVzA5vvfkRKf+SCW9L2wM67AFnSbVaEiSYqYf3wIT/3dGByEhGc4SURVdDZJ/J7LLfefzMzLK
7ZgqTsN2oO6UK/+d2fqXAPQEdLh2Kft0BCF3kfDJpPazh94IbAc8aUYvo3AWEcCTbMUr3RAQ/CZ8
yY03XYYcv5E5eiDQjpVyKMz6yOp6SXbZvpSVUSMaFI8F/w1NKGRWZK4C6RqoDhw24A6ZSwGbDm6N
ISEhLcJNe67jS19GD0HoZkCj+nKc7O2ki/h498NwDuhMNkEUyJPMW4VwSDKWAIKY9VOQ6n+C3+dG
h5bzrAn4yXVljSKjbcZd0b1jAuhQsnRhD9KsDIcmjFldIljncdSduvGZbZKQj8+Ior+3RfDuRTTt
J0MYvvqWiR7+8PVuEDfY5YmSs3t1JXxSzxuF0xkJ3e6aEEngG38bejXp5kt8ZaVUsZNniuZla2Qe
0opNDBvcN3zzEW8FX5n+xvuIYzG3CChafJnaztzDmq3NPdxvLKxVONZOmo+2aCakWGufD53YVZSp
l5aN7HMKwawHUmWG4oFibWyUlUJAtIGmIAiDQgebP91ab9gdwRsMA8RURx/eqRB/WFo7hgBTmBm3
r/s5YCGaN/l+rU+fKZ8jn0Wkvqgr68/ZxI5JpVHWboct+I9JdshiVD+0BFJBdPz1VFtAsSU5VDvh
SUzVbSrHOT9ccPeT0bJ6x5rBCwidR/D8uFxm+jbJgCXMj+bgl3CoLlTe8/YNM+9H/YWfULs9Jq3r
xlBQLyB+N72O29AyTejQcfCW2Irb7U4tK+lRQBb1sXlklooDrEuJmdXwQQcJwWEyFPgkZM4ET0ak
/RTwmAh66BZuK52a6AF8H+GYuvpwooOWGGe4o7pYfKy8vayy8MHDv0L48J2hnIyEbFuSNxKP5Hr1
z7X9ViRko4EIHXGioI2XZGM7zy2x3fQnoxu0mTv2+jgZhXgiMf/M9/8YspI2ATLiyWstb4b7SbUX
iHxSWWuyH7TG12R748mWe+TjeNPhGG58vdl4XoZvplvYjvEQR+7AnQzsR2rW0HxUwyVQGikYFs22
pTL2YpJHxsNPlRSiQjvpEcgmRJCzyJkg06JM0XnQ5S0rDKN4P5VULgGBEWezHEjPks4HsdRGIEB+
ZPeOynMYezjwC2BDjkV9AItLf1blsaJnj2bWtdOR/GWIrN1wz896PaqPfYzM21pGJOjC5HqOQpTn
BdczYK4yUzzpDuYTKhoWP0fSsoxG1CKY3Rxx22RAle2vll6M+NytlqwytniDBxH+i9Lbw99NzTvG
bMrJlnnrw4FGHypfiVGrt4xaL2MtDeQAxIUqeqtWCWbKxqSmj24gYWNRZIn8M7qNQe4fOBwe+59p
5EvFaYQqjsHyuJTHvwoZrb9ztS4eTC9ELchYDkHPNTmxmcLMh5dNtKnhdZiVJiQiWnwhlv98HeFx
RsnaHj1SvvcR/jOBHLy0GviKS9OrjTyYO7QmK8KlVYTnw4JfksIwcB/uWcEewdNUrjchyDPso+oB
YBikAo93gdggKSD3FfQZ5j+ZPpWP5UgdoKhd7ouAGUZ4LjDv7mU6CZULwNimrN8eaXywxdKfLlNu
LEqmWY5t0006Qsr6n+PpszmNkn3uWQolb0ipOd/vaN+q4k/jtpIShz8cVioLAkFJGSN/n3f9nJH1
EKnuox21ThhV0UCrTFpwKONLt3SzYQbu9nXRcmG2soKAJXypqPKC0tcLKUaQy7peKCRwPRK6O5Ps
3rkSSkdImM+59s5krjv9Z4E7wTXxYXPMAf4fgWlA7vHXMKY5TWiAkc53RoGVQQd0zxycywhg4z/N
jmeF9TvmJeAcyNW9uOEBnZeWaRVTWvSFw7tfYld75a1c07f7D76V+2DXZ0dHDx4j1EsNJWszN8+5
4EWLsE6GkCzrBkYVZtwf1xbMbCgsh4TfVhRYFfXWp4rXsjHtcM5hvAdTusaPE01BEaDWGwu5Ob3I
xF4Ql47Vo4oiXlL52ET++mjEb77rBD86k1l5aafnrjrsqw6jeGPnBeV8cwVxy6sRvXhauB+WALZQ
nwKHCzmKWOZ5tN5m/NDhxwHVcuLlNacTfOolvWP3jnXHBuPWEB84UZGM0JZRusBkeW8YNgDpxB8R
SkDQC215yhohHKYdb0QsXF5RGauofFmYLeA5bRLEhTsDJfUgfXx2s9sArat8rOu+GoOG9+7ycE6Z
q2hVr+Rb31i9szLugkr0YBvuve7BQNRPAyiH8q/f62fGpOuzQSGujy4NwEaYsELJbv1d0/C2Yg8E
2vAjQVZ6f4dm2eli6tYb0sHEjaaQUejfcWTugn5Ha5Tk2WJLP/KT4GfJgzqkNIuoIlmQ0g8isrl3
wukTWl84yo12m40KlvMLEUenPQ46Rq82iIYhIZYbSS5z76yz3d6yWfD4Y0/itaUbrJ6gaXv24GMU
elOIHkBr3AE8w9cNtCIzC2HArwraF1TGCErs8ylQHG/Y26xdWcCz9z/59Yz1GaN/iKehcJwVRwgt
LMunp6bUOd0YIEJXHCv1WDOpu/pW0kEjjaAqU/wxGQ0PqFA3TFDk2dxnGZ6tGdHSpCWiDkf98nLm
IIOBe2SWpyhaAP+735TgjrDZm6CXNiMUbn8Jy/NUneE0UxSJ7JRLBv1mJ0BfqMXV0u+THrdK5f22
ZlzttsIL+O52VSnupCSGtfJv1XVj7wW+AkNYyvSLFdrb41v4SiBNOrN/eWrwz0Y9lsDttZAYk9Ym
rejCJ4slMpBt2jeAGctzARmbrNswQlb+PVO0+W3+beuR3XSky2oNYfU/BDLv/kuSIE4H3yGgiaqd
PCBKOwt0P1t7tpBdyd+I0FSGQSFlvglKXn3nJSTtjYEhRD0MqFQkxCGfIhfXVAUtnd/o+4yMCBJk
ZSpcRYlCNerzJ5Wko5nGtyaWmNBJV/FV2e6uPNkYzVm+GKOqMf3lP3u2UH5K6YHW87QAM/jUuf/y
mS3lH4JQbDWAhLfnh7OxMH22l5i6tVWOVa9JSKz0bXmmBrdwTUqO0IRcyZrQwRUbLT/wuwnTiKCi
ZTffwFuKaglfweQTU809QizfKO937FHlgAyffcrnt+HMk27DKBmEai0t2InZwOfImLEsH4HgaEA1
3PBh+nzZmjeM+Wu8ld7JqePj1BdvjM7/bTUePiauiGunXMVlezOeFZxSeYO2gEW86QxlYUG4ASne
88+5UhDkgvu+f/x14/4E11OcRY1Agaod7Eo3JC5qrCvRaeJ2CacZaP5llmayX7ED9If0BAALr1S/
NeJPPemn4PuQUoXThCdyWlhLTxI8UDVKDl7m6kEgDodFQeoJE4QluLhwDk851EvdvZMFIDIFTtgt
0CtJhzobM7cCbQpWcGr4ARhksQD8K2NDpoyZM6CmZ2psm7U5DvrnuH5rvE0X3jHXQsd3l4fKXKBK
KrGMl0acxxF+HZ+fMwJf3QbYXdiaIPp9AWNR9QQ0fh2FFAcf1+nCRotcTNMERppOI1YDn8WgotA6
z3mybsVJ+mOYZfElNevh65IMJdEBT18gBp6TBmFcZ8NuEqNtLW5sZ2xX7huGUpbPY2dU+xUMZeES
pFv92z6YU0J0KGDTiu3rjH60uYFSmHoiiPlTDOa6Qco3XCb9wGugIezxSa0ceSUq/m1Zsf8o9FkR
Jqlqmx+pAEsq4mTmrGM8qx/QTytbCo+I7iO0rGZrLQLli9n83ClK8oDvu25Cjlzss/r754hczDKO
BRTeuyyHtdF1Q+683i5j7D30eELFXcRBwfDmlkPgog1m1iWYg6D/vVlV33sIWRDtN0tZcv37gUkq
n86/URA8bMPV+m4TX7GZH3NkR1RREAVvwwVsUcOcIPc7K52Tn7paJcKuUIfPgYIhmIxw+ZhZz17w
Wg5INNnAaYJZtgDnfE4asiOiwMaip1ZClCY/F3T3WBsrb0JvVW0pCv38GtYpCul/Ov5WDpGBezHX
sUXyVou9zjZxIAQRFN2zzayd73UdEPLJIHcoGtdVplQOVlzvNbOTf9rzYLRUtz4kDdgVsf1YJfSP
RgjC+IbC2GcoO5MASR8khLdQJe3CIs2blm/O+OQr4r6uQ2DrkimTK6sSvjKTD7FW73/hIEXd1GE+
w4wnCuIEhsEWCv2441MiLTF5oyJEbXQfcotmD52INS1yZYxfrC9v6V1uCjMa6Lu1b0mWFqJNCFuk
e0BqL9sL10Qxidsd9EKEe+QIjw/nP7LX65TYJ8Rifjw3HyXOI1JonmB73xVqAgSOVmR/VrLzgA59
H947vc4Yt45WeLmynHA94oiO8xgw52r4addteh2ZPK+Jms1J5kbrHZPLgGYU2KCaw+7fyA9gBkfO
Tg4n0FWw/ZRJrbrXtLjiOdOA1W449X1w3Xk/YDJEnLHXPHSDcOgAto/Ch+ZIlQFn5DjCk3wzqcEO
EOxn66ZARbyJOOLh8URJIL1WxyuT/dLpK2Q4vJ2x3eOvpJHjP81MmN0Y217KPXQqi8mUh4O9CK5h
kjwO9SIcrgPwQwQXZBrlWwvBfqxoNuKYXS2gAs/A4/71O7xlEbuyPBsyyZoqSeSrDvnED6LX+uiw
E6ld9oRLNWTxXBdPH/E4zzMiRmNuqkW3bPF29XA5HszUE9NKfEEhEAb7V0fVnPtkit0Vg7mT4ZQG
mE3MTbZocO8VPMkTxxxRBzap8kyxPlA3ZmFe47ByS/wwRDTs5VpkThbUufGhjDEt8Sb1DUToHams
Y9/IIjvU8/eOOWyfZal3LkFnAMkekBJ6NvIJKmqLGENnikhV5Kvk8+tBvuWN76y8inXRf1ygrnha
tZTb0DApYCQA7PmYDgWLM11avXwPpqrkH66JI6xlAT8a8i7RExvSnjoTgpzS8NrVnk4+E6M3wwiE
8D0/vr1p2sTvHVbAP4HrTkzNUD5GRwox4CKqxI3BjUvNnqyTFQNNNUdoVo/o2kyifhApwrXDTFpM
qwAKMCFxrXplXSk8fXr+x1Jm3nwrjhFCPyplUmCqHv5yU36SEY5R6W7tpBrTGgwF0hR+9sVMN3qs
3m8uEb2gHeRG3qVhRL5e40resR5rJeVw9rHEY4r0+UL+6iANMJG9q4n9B1BlNdOnxEeOKSLb7KG7
GoCJ31XA0QvlPCxcZddbnZrd8v5gZbJGqwIGDjjhU1bFyJURQm3CDGDSjKBSRcZF2bbqtaKxg7O9
I/gVFB1TxMLSqpQ2u6svTihuA9RJ99nVfhvSCz2wzz5EIV9WrpepM+XRqxUwQEK6q7m/4BPmVdM+
nhk6HpTm3NFUwOf4qB+uITTScxqfNl/K3JrWSQJE7KDaBBK1kZR3QrLAB4jCPiUgHEQ1koXd62r8
olXe7fwrZNCSGKMwQStkc2UVCDR45H6ocyd2NTeyLcXqFNVsGMU2cK3s7A/hXWUe5cipQyLYVFJm
9Z/WbkWcazkAYvbhtEmFrhEpnyXm37RVvgQ4tXb3914JN3jtNbvb9kdjpnIEE4T4uxI8ipl5Xh51
ovtSj9zrQHAMtX1f6a21qWR7GYv5DqxrwkOS9SIKbYjAHzgb+4LbV9rO4sX1gZZdzxt+uSKAM6Oi
R6EiWd++T3HR3mkSXjr7jh8O29XYk/0JL45Dx3pMlpTbseQY+MhuvI/jnIfl4zzkSJx6m33wXFlj
fB/GtNCo3BdeoxgsI/+Vs5y4C/ZB1hFOlwQvnh1seGnop7imhGDMcaY6CMgzVvs59V0i6qqpE4Rg
aCMN1okLV8RMncgskSdOKTISCLGULD58hj4zHO42/Vs7nruTOT0VsXbbGmSEa2EMpJ6B5HYCVCMK
pz0K0g+3l27g5ugWTs/ThlQPK/qY1sybHYKsyjSVOHW6cWSiRveTQHPzexld4t2KX/jc0ZktmAbY
iYGVOT9dK4Xpn4ftXvvmge0xQUtdDHrwIskH0riSZM1qAt2cV3OtEPBqVs04Oem0k7vtS1pXBL25
OQkR5ruTzu+2X7FX6q5rcThCVAT3pteDH/ZmHqFtuNSe9cTBk/G9lVoikKGgXvNaXRk6r5OrXsTN
Su9t17vaWC9d+z0WjO6GWophcYCaCZ0CBOpp/qG3uJp/nuhqcRHIK72NCsmGRT3h+ptr4j3upDY6
x/fgyL7kNG2ZOjzbu8HBXzyliJVTF27azlHXcClA5Gs3U4Y4hVAlsxMwepvQenGXrZ2t7qx0IcUx
delkWPUcdHI5PyrLFZNHr2pyNBAaHZ1GS6yQUlJnGd7EkRIn8N1icXgNtspyKhoPt1cNaYENrXr3
Mk104uyIPE0cSSs+mfitaYxStmlCmt2hVRjDs+7El2Tf/lyklA36qcVDofuRMi+2pT+ENyWDeiGO
sAbYZY6zYn3LFI3mQkyQZ70//LtgUNqy0dRorboG611OU2ICbdnmGQWkt2m0ljhHOSzPt9odyKpZ
RO79lkSvaghGdLrVruqxOLg5DbEWm+sXdV9lbgEg43yt86ouDbjyN2hCnMyon9pH06hSd87tNggl
cgEExQ1/p2ViakkYzW/70sIy5oJMQXm1bF1c0+taKjm5Xi6LPCvwmDBvF5TYjEqfuyy8FHX9TA7H
a4z7y8Vl1cAp/DxQJdo+saU0A0fc8N2PjGo1Tf1nJpnOKlPL0P07A81jUKrTJ8Uvdagz9VmaY8ce
eS5PULQmu8qw7kuWyGLS0jsZ9lzcQPRNo+9sILu4ShGBeFCs9PwV5j99MWE9slWCYhPLoXypGKZo
t/sXsAvC7bPYXm0hfY08UW7j74metB8LyMATgDEfn4R/20EskENXIIVyb9KDJ1zlibtfH+vhyt6c
NsevYMbvJ2S8VDO/WbvO/Ugb335uQSeSGFN6KPNBERjX29LRwQ9w/OSGkQrCJlfRZXvAwZ1ofAgc
jklHz+5MSh58xnAeUJL/nnXLWGgNFnq1NbANcfQwvAjX4HIVZr9MklYf/so7MuYQVIqVhLTwWgOV
HlNhx5xWsYE9evDkRUePZ7fM8IrQ3eB2Vwqnv02ahNa3ZU9/JLhEUelshxcRVYBvyZpSgu4rHYwo
pMAmuNvxumLwpRb2WkbT/M3B+fR9Hy3a/oHanMTevgqVkbOz8AWg68EML+odM6Nivi9nXpwY8bqh
aueO71FvVpOl4eVXV8KXGfYIMatYEPsLQUezvYWEy3NjCrPJwH1nbTIOsiTOT/+IF7uikn6ei4oY
Vy0dpFiVtR+pyH3p62/as0FTKRRUkEW9LcKRqtx4E8n9sDfVNjLxjktOiVCRLmCpf1hCQHDIj8pJ
R6488LGMjKJLH8f2QGXVVPr2s1/sV375yQa8boZJYnX0vHpKHT4wKzrvmuVTzPFREb5wu6xJZ5Mu
o39FnQy8HpTgkVySe9nRaJS0sU0Nf3wl8gWaAc9RSp5JqElpbE7uQHjxsFgUSheDFORl/LcAoWPL
9RPadce+Z3dkNmGsuhmdDmO80JbMAYEYfZbqkxsw6zaUuLmpe4UdC+lWPkEseIKTHoyOg+phfnyh
YMrWLyvkjIxYBAoe57EU7KyPPBtVdJ8ScvCwH3hzNbxXW/wOiaZ/oR5fYRk5dNrkCde+clzgAtSw
daxxwbKjWyg2mCvIz2O/+a5dcurCkg3EEtCJtAMHFyYpe4jk0Soqq6QkwEFOBMM/hkQIQMn9iPZ+
jxzFnZ1DYvsCHykUg+fnyYHawIxwpN8lsaHc7t6xufE+eZDuav66ErByRHWrouxFEUsnEKbBQN6y
noxhY6CTGXyBX44cxtjDh0ygSqTYiuPn9wEbRaLtMsVKSZ4iMI3WcjfBw8GM/2WADxAEQ/Sc+RWu
DN3Ro0SVpVRZgT/ThkUDP1vE3gFR6MoEmEl/OKVapyr9XYJ/sMhNjmDym/f5VOf4gYPrNWPlLRZp
Q0Ws+iM2t6m/2EA1SYZeja/P5aag6kO/JmJNxci7wDURrueK3OkNfs60weEVBIhUysYlC40rwsCd
7/v4oTpHd16X1JkqEDWqM7WLRYY78n6cbmzeZF+PDC0wZlbNmQJXYG2EJwLcEE6MIB5jS5ZIjwm3
bpGXyf/jZ5mQx1dX8m22J76vqYw08PI7uQFnKTky5XsCAcelnbiRenybru74FIsQVxsGiXWVYpIL
0y3agTrZGj+loN8is+MPP3na8Xl1gdFQfeu8mz9FALR8Cef5JPib1cHTPKdpSftPYdhBbIi1eNqU
PY22SdMRjVUGEs5u+otk+GicpSiEmBwE5ItH0W/Ejkveoo4vHDiAYhICPHIt4mO5/Xv6aiD++Df6
kaKScNZYzYMYCCRbXouMIR7L4bSbDjuMOi6LWiZr4kdahUSl2H60OQbXL2s7YpQrThm5DQDoNnLE
pPMND+FVvAzD/69w5nR/lnl4n12pfrD4igaOYhv+S8qF+YNt6iceLiVg3nIQfDpOQQVSX3eZ7LEn
9PLP2zkaoO5eScXcs6h4aveKLPn46uHDwVg/fK2uVh778674scp/ZVxSdv8VUl94dK4z+r112zOL
6YJaFKqdf6ggCW3L/vTAiC2iuxd/C7jxexBXz37tabF9FZj90KQAGlKcflZVaXah2w+EIsLCeHp2
mSRvdzrnOeScBRoq2T/jljJnniHpBnWmBSvuwPsy0nvQYm3NodHE1F31987Ek6MvINoimyDRtnYa
gVH9UunlWWUf8OxljpMnxcKxUcrUtt25A811AuXuBCApQe3a3rwgqPhVHiQCZcIa4KPGwNRZ365m
KFZxJpyBIsWCL0/4V1HS6r5QHOsGrVDpiEeZQR9yibE5tldh1e3CDFL7hwT3wPQInz1ihpa8pQ9g
JhxfxJridlW/fKnEvWZJQIlDmbfxnVvgl3zbkCMZTBYObinseNZRHN9qIR14FjvSDz6BeWcUP4Qq
EO1uaxTzYQHZ0hLibbLAW0/pzLrMuwnSVJJrf2NUEDi+/moIbr7xk6GP5dCAt70QVPLqIkVZ1qDD
U08zbxrZytz9/85dwbNF6WXyAs+H7N59LLVDB1M5fX4U7FpRtysTA4tsYBGcayJ+Mik1oSuMkjMU
SbcwGUSd/dUojFwquDwaFsSm8jTQv5QLV3l1CfwqmzHyiVgy2zxB397v/TWybFTcZpQk6rQoE9m4
W/RTseiwkGUQaPe97SCTdB2NDL9jOtFxFtVVRi6dRSr7HH+WRVgN/uGmJcvOfE7QwOFCa8AuRDjK
g2/vsDtQ7eOhm92BwiMb8Oqv70TzgbSer5IxKsOVJ6xq6iMl6tPIDIFaf3Krbhkrw9d7UlYRqp/h
49hmTN16uyJqYUpvMDv9vLTHuFZ4HXPtpAXTd1+HPamZDZ4bKO+F9L1VvUmZPnjL6DamjO95oI7w
kha/BDdrMels86/y605vZWZpkXn4SZJEr0HWjqIa8PVQXr+T376oo/dsUftSd30fL1NF26OCP8+2
tr4ZvF8f7glo7Icm+YO2es3r2zQUg6ngTn33A7H0HyseqZSN5ReUQiGJ9WdZmEG4qNHyTX0LkIPT
6TSnAiUC0VkNuZ/2a590q1sUEILhyiLpU8GztFuUTlhMGtganr8TBcGGi4/x9x+x9/JNd+bIQpFq
kTnGgh/FQu41PxfpzLBlDHtFjiLWpP/DTJ8B1h93SEIQqAxkghBLQUqCliAKHLtvFGllXBYFkzJF
yzuMKLdXmStq8g6Vg+DeDOJV1yMqcXfVS5in5FQYZ2s271EPRs3qZjX5oQeGb+Z5+xlTY4IKu2G6
nLFKHDMVKPZH5xzmkY2TiqBlvtYttU8AmH26r6gp/sygJHl7Vv+yOZ7Yj+jNVk82ZvEY14kNiGEI
FP8S0ZQJRT6xIBfWrQQROE6tyxSczmRQO0VH5Yb/4r7mMoZPtl0VFfaeUhZrgFEcFyQbLSrwV0dK
anv1MPaMheYJPV7hkp9RqhCIsH22E9CJ+lLBUUYAd+JvJ8USQPYid/Td1XYffS5SPp/5DzPV3zF6
Qqh8+JGid6mvpxmk65/hBedoivQ540lIDZarPRxWhzfHj+TWSwy83cJGRpDdib695wnhz9Js96Wt
vum9ZF7lTkGkvLtTSUVnoKzTlAGUP50RwM0Fc8L/5Ji/iNXfN/JCmtCDpoFV0N9im36OJKGlBIFQ
TrqIFjeoeSYAbJ5jBsrBNXbdEkWnmtrCkBBC9+X/4AGUnRGALeOIvp9FHaNdPzgPfnKgxCyH4Ra6
Bot1RvftlfSGaTwM6K5DaMPIdSbpB2YIKWB5dSH0MoRyUXvNyhRhi3o3flGlYTF6dtZ3kHo/KbtV
7jNJ1AVz1uXNiW7R7PMYmKosVihhwbUQcD0Y7PEcjlyHJgrXU6Bhz8w5nSRlBp/glt39s2z9qK9V
AiXqDpmUvL/VqIMublYjVxnrlwDCiDxaBA9sTIQQayJbaP3bcvhmaRiTirOgOU1kDw4A/lDYaEvn
xty4TgcvaQtR5tC3FnON6jxOZwyr9xCwzbHMoAaeK7E6CG/JXwCfMj922iWrqr6ecGJzPniLv0OA
Lc5irZM0TaMxKg0aivPg91b6ny6V/Vk34ACr5xn2DC2KXQlZmISPA2Qlyy7FtMwXPM4EXeLnaOzh
e1wWkoRz/6mMtsz0Hq/GTUOwtp+8HEAfDzhn0fFC4z82h6QyJA0iPN7YmPsBMbHEHTqR9+Dkr5nX
G80dvmMgYyLZ7p6zDcTLHZdnKX9ZZaT4a/2dYtbt22BGCSAE5LEGOeCJmU4SnDHeDkkVzUSOKp8d
9xW7C5Z/tKexdmdzYvfTh6vFXWai4LKNokIHoeluPjn6zB1jWLScCWEAulLuPXJxzHJkeIkN+k27
eL8KEeh8YAXGTVUMjG2vfsdgSxcts6CWexEK3kS1Ac8RU28W1a5N3xtzyVMjT6M1LcmBpsTJiUuO
ZQRufz5JqzQD+HRvBh12VVszAxPWRDvNmhjDCdSBq/oxzFlCdJJb1ZUmJwFXhhZZoL4ZEatwNIq/
U+fEnJxzWIgM+IVVneTgaPvnFiodKDFiD7LC8fGeUxYziEgz0bL3oOWCQ7cNbcnyy6/Eph5ktnJe
UsvTVa1yzXiIIUpUuZ3fcAPp6UvgWI0aXhDySmIa8DJCDJcDGIT6JDfHpOeZTh2C7WMOQDJk7YOk
Cd0vaTcsTixp9M9ghx6dHQM21K+cHdZ0fd0NnLVn9hkoYPLG+E+3Qz128V6iBWx+2mOzVoi50kxn
hoWEJurgmvgojyYiDfitpmswMzUNmhFWV3N7bo16ux0UnQawSULuIZ5Y1S70lu2fBjBTNbGiNCkS
61cY0pw0EX3nv8z78oD6UsiwAlspoKXv9MMY4GuRCMQN3zXSIIC/fSOVZzclvzFyj7CC8iYzdWTL
EADEgYAf+Vq0Tp8QXLTgi402lFgUmmrMac+3MXmWxRllS+8RZKI3AZW+VDLkZf+V5CXOmWjlIXOx
GWc4tHVI13uznKNJfFyXSglj1dORL2NAgbOcQJf4IJ6B1RL8PgOqqx8+PWwJIa0xjyFlXJmtXXx8
XDmGSwAiKwZFvUNLPWpEhm7rLC8NOVYBj2XxTrq/bcGhhK/2HzXZHtyVHC1PKk5P7rExMsK2xfoB
5pAJGDoRpumNVt7CKyxsyZkAPOv+z+MdfCHAH8HjVaKT5AAfX3qCDv/yPq4blhy9HWRzDzYi4I7X
qcN6wiA5H/IXcdyRPrF7phmwrFdoGzZT2vNFKE+fnymX3tYyVyS01Sx5QhPvzG1iWxuzO5IcQm1/
NgWX/QEqe7GX8XtRMPOh65IAe42Lg1MJ9yVxNc5U9SslFOioxeBV6+N6bkslbhqPzhYFfzz99Jxy
TeGhCD6zt3TIbjVJl6FIbqhn2Ltvo14Dj4a9Lzuouj1LZ+VFPUCtyLa/twjgmvbCxrdnvPeMMxgx
XTKCA9leTfFJbrfn/tMCs/d97SyLQvCI3YAJWoAdNp8aCpmkUCiNbX6CvFN1e0NOKtfWPsoyDzNQ
WlgdNhwNZ5WtCi2ebKCmZQu2cM1GLId/3asFoa732EtlJCP2eTSAmZWIKRtrw9DG++nNOIiFMATa
fOoqufsv7ZoX4r4dSI/xan/LkRub2rvRaLv3ePQhuoG3bIYy0PIN3FDt70JvH0M6hTx5ieiIkdB5
MzDMtf/T9ZmazxinsjYiCzLitbdxCSd5Xp9X7nQG98PEhZK4YbG8NYEECI4w8lVZciLpS+a0rvDu
CPTkvMLRvr4Pcwx97SPyXhzSbDfyXrqEi6vkt7oDOFjcPpbiZQQtM1/VdKW98B/dV8jUGpk+gMPT
VoRI1wPEytQ75PYr3xV0uCR+KLdP26MQXGign6b8YbuzdQq8p0X+FW8Qxj49xdALqrIv9ymB7WBL
SdnJRosEMSi7NYKGjXXMhR5jjmsB+U5QQhU/pxADS23bcxVMOPM3aGQLZtMaGba5WFAe0g6tvan8
o9ezaV3vDDmIZD0+H25SkUViYfLiIOA3xsL5DYyq5fYxdL5SYCESC+c/cDz4IKnIccxBjeoS3D2A
Z2ITKwmrxiH11I1a9mlkTmVvxysVeg2h+V7nz117q7MUY3Djn7mzZnXdK06dyAjBH7kLUkjAWlmT
419a2Y//gMWCOL437TKbsl21kuTGCC36OJihHq7Q/BuYPQf4oqahOtdquITLtfangkrUQ+VuWQo2
Omtlv+YgPEu54hAhnYG1DzdFqBj0+KPmyaz/zP1Vwmm23W+q1Ev4QvG9rA7pbbK2MUFJN3Y6SO8c
2z+ZONwOJXpCI6VsGxiklstRV3zmxcDZl9jbiauP9X6eTSNfs01fBPANGdwTQWU8rnzCbtkT176N
FZqehDnuwTs8RwIR4FQfR16/LBZuapBYeDeWdekh4D6o/BdfMBWt+nz1Ww8z62dMrapBjpXYaX+I
Gbf07Ke0fqO+A0r9HMlyqD0wkGcqg8iVHADGV/FMU4O29ZhRvGL3fDgalWGKbqe8MMHoI2dWOkzr
sMVGqnWH8gAT2hKCUVA/B24JgKYZ3wvaH94bYNPEXeIwsig6aYGMq1uh4FNKd0IqTJYbiwZnyMG7
TRqVu1XKX8SJrKTUAmGQxYb6ETcswoMIyZSg7MWwUcrwvqS6PfvhYbfvOjNxK7vkOQPXnHZfpq61
sGFi4XqKVoOMq9KQ1a0gZlDoFrBk7kUiz4LfZolMqYhNWyzPbtj8Td/DD4HYmKtdbhKvz69jeu4w
U4aHfY2jG59VGsdzLT7PXmTTK6zPXOxO5N/AUxnPsCpaIv0hAh2vPJ3PC9MjefjmooqJoBu3qaOC
ZDL4xXl3jJg9Oq0534qjL/v4wUt+CF9ndb18MFwd5nTAIWphvHj62Mv7rBPuEkC4yTH8nRkXW4gY
Fa8+rusPh0l3fRh/JhNlCnbg6B8/kUdxmPIrCxQkR4FtDdIwwYA0jEOliSElPNwn+TGIhHivHijo
c1AULoPhDCP58cnAMsl+9ra4UQFgjT/n/9vxrNHN11YUEhXTZiZUruOOhafvK4lw2IM5Zp/fB6mg
oZog/o9DbTOCGxYvtfr2jMNynDTPueQr4dpCSxcgvKN8quSYlVMIRBAszgQDHzu5nHreIBX3kE8e
cW8HrbOW/Swp8oDlDY5NrpRK0vYbZSXznARooCq2CLS4ItEXxp4CFTkyejtiZDNUlqA/AShApv4j
UKgBYBemxirxYVGH3mrpEGfVl9BQaTlKEEiC9Twq7NWDXCiZDfHwjrjQe87WIhbmPJfZpnMM9Ta7
0Gcf9ZedpRmDiUpsXqInYOlaFF8AEXgc2KOYpn5gglU8rSXROkKM1QvKxrofIVDiyH+7RVExTul7
v9huZFJm9nlT0RxZMfchD2bZhNqVgwnsJMTTcicrOQXus9guN5ZPK3OXazfNIa5GNiU9Ee0mFvtx
bCq+rnvLCwi4Fqks9QN/r9sqdM7+bWTEmVmqOsFoHgYMLRoZh8MXHfONgUYAzkR6iGKZpsxYvCT8
onZSokJMraY/qNvuc3FGdZ1EER/LC+5YL6sXnEwLUdYjbLh7HvsxfMZmun+biiDZlEGCfclTGNiU
Ge1inTTaDLcixNZHVTmmdoOa8ojWJJoxm5/+pyjk55Pinlo3KbOi2CbIuTElejhpmh0AaBvbXZ8N
UEHaUyWFajdkoVS6aJYbUAZDDQrYiaYhYw0VK+YL7TyGtXJWgkQJbvMuMDzJ21HWBnwKqbxjuk1R
APu/6/mC3HwZHYqRsDZ6qcdNg5yOyw6LZCrz1mfC4EQ8fTSEBibEpNg6CpWYxlnQr+cdoY81b91+
rmfSaTI1MZ5x1pKHKNVU7XOJmjlyx5ZTAC5T/fxdmsvTLeFcpcBFjwAlZiNSUgYn64mChKRo44Aj
vbFubRVGVm3HCWN7l+jBBctMvP8zYnjDbllCIDdrdDvTqAvc4IM6/Kbazc8lvbzUWtPhOJk6rTqV
9qcSM6tuDFZ4qzUY+ZPKmO8p3vNTsxjI7fMbTIrelizemcQshUSdmSJX/PpPGWdJz3yaQSjhGK5i
3feq/XnOapPo/STTuUVLFPNVBhGLvybL7hUWMyygNYRLrKS5q+0D2rTv0u/xHDbi2JV5Zx9ds7Qm
wz2phzhS7cKfmTna7WlYsJfLsqRV/1vfQ5IDPASsmgL1EG0dSg44/ZXdhHWuSXclntX2FrTpflM8
UWSoTLyD7vuXiIbtshmSuaa6rncYAVFF+HhWoTAGPsy3aG9ZvqcjuZuPpV0QT+3A/5A5gEjq4rBH
HfGdh6sPWMyDltI/s1hB1oppdxq6PLfnh8s/QZrWH9ymvYyJ9GWqrrW/s+nHVeF7G18KRYUpT785
3FFcawUSLci25lUocArooKOUacL9GwvxXP4sMxXjEFkn1lZG49cRZWuTINX3P6Zq2EToxPuJv0x+
MgBc0lse1xsYdFylzFXRKP8ysGlwig9DNhHov8UuCbiPvpMDDVtPxamyPG4tF0oHmF+qZ92Mao2C
U/rRBQa35/j5KRVIqp4FQhShT6dxEzrlNnUweOos5nO1zc1i6wotc3z4TmwWSp9CtO+R1ZtGwEVl
XXdVxhbbtRi8EsQekttaOratlTmXUZ/PowF+3MRIyg3OHy5I2zImbgqv658Nu82eca8F1ah5w/Zo
ppcHKkTKXIvgieRuXDtpaNHTCSyJE1ODB/+JEyj640nvLRCFYCdVKh4H2EwJBZNTRwl2CF3B0kBO
GUe+g9GR8jvxDujWbq1nYxOeJZ3Q1z7ntgabv8UzBTDEhdduYTcwdE1NJZ6thFjSBeZC3ORkDl6E
TAu2ca6bM9f9xBsySh/emU6VWZiUV/KiuUmxtwSBy5peoS3dz830xLDJ33VeyBR1fJtP5UysztVV
mBXU6JiIgx9DyvG7UQsXK2UPDo+0h47NGWoW4t+YIxPhJ32gsR+UqBuvjOqjm4t1YBMVGQdtXSAi
8qvn5xIRFjhBzyPT2IgV3ehwbrLn7Dzj3rvwQ+roEvUujrUS0JT8IxUp/ncibKOhzqexOxbXOc59
RfkCPmwDK9WV3/vQQnSm49BCOB/SKUHF9v/DdtIpvhMe+JLHzzEl+cwAQJkJpC5UO14zsy0OI7Vb
YPvfk5+48V1r0uns5y0csokfBJRA5enayheCtiYSf1u2mjCZ1eEPpCr7Di7wbtLOxtuqJl2bk2j7
ZbIgcFV+9TXqIMYWAWD6IkIj8tunGnjNKgTDocBrqeuQ5ppnlwh1QQnnYkH/BDmf4ud1Cot2ChCn
Kjr+6lLh9bS5PrzocvGdkJDthLMpWf4Hh1IpvSSY82q0ZepPyy8qqjAm7IaSw2YCdhf9COq8NMP+
w5SlhfefClnpv2oOMf+wWMn5Ax9sZDikwGz+haZ+lNk+dwODt9WFzxSzfOAhljVL0sFtpEbXm6Dw
ewNFZpdG+u5vy8I5DZ+724HCnFnQNePIFfBLgU9C4rq99Ydrp1YkFKiosei7asTawyfn7wKx8Cms
xZvTkfgH2BXxm5nqoPe15/yVOVzBChRPuLc/kT0DilTSYfQLbgk9Wq3NP6MrFhNXCETQn19lCDLh
ISFe03TGFWzAoMSI23uHo0irKTO3yjcOXwOgd/fvEjPfr0EYYbQ6ORm3KXBCJ/wlXg0prKuPEZ4i
cso9nEA1vjHThUgO/+c4F9KqlK2tAQNdDRQ2nR9PJrSDKLjYdH78pojZUKy54vs0/SdnB+c0q/lg
orOfpCnSJGaorObwcD+aN7sFdrnT66VHG6go30aHPF7sTP9i179Hi4rcOs5CaxyMDRIIuyDbrsZf
d5djzwPL6lihYbmZwi/Br2rkjr7plTmTq1lTKjtOtSDArgurpXUt4Ume18r3k1nmkauEVZPaZe9F
q7E9p+OeaqkKukTFHH3n9xOFFzBUT7WAg5UaogRMOaW7IXjApLp0fJF/wae5PU5zUXPfdwuVuFWs
lEY0+4mE3k8mqnDxiYKkpJLcuQYfRfkcCMNR1frorRMV+OpFhC9Uu75XJNksaLy09NgDMKG2OyaX
A1xJ9D7i1MV4n/8mQUxVNIiPqqvA0QlyA/4gBGE2J1AlZsOPh24lx2wpt3lqP1n3fZ/5W4yiV9VB
KFt0Wzkl1fr4EBN42NBkBgNGmjukdqiBOZBIHmzYaSXc8rAp+tB+bJtcZVYZTct2nRRrFmUPI45K
dMb1cMObfIVd/k3Zt/fZJoRctSN6FLZ04zSKKv8aKB9c6toSdddZVUIUVCP53adaOzc1lc5+vVed
TO6nKM71MHY0nsQpT1bNMfqkmdFRbRdm+75ZLq7a6tVqHoMiyUJNp9DPl7UdwHMX4a79on5JPf2R
ZL9PUvups5Yxc5FvhprFJXuuwLhYtFsvmRKRFEOJuRSV5y0p8ABNe0BNKIVepPK42XHQTRxyr4z4
4QXjLSMxtCXzGWUvDE6q1lvlXo0JI4jCTS9xDiXjJpldb4t5MiiwThvTuyN9+uJWPAvzDV/vvHpL
CUyrc3Kz8JwU0ZHGAORcVJFt9srsrGkLbzAIA/HLSnQkYQdviCF95LAyhpkwAW/jjbkaKO380pOm
aZQmhhDk2EaP8NP1kaP1J7LgzFF3VfNjOXMK9n2TVlEZxk+af7z4Gf3Zob/+W/G6cfhaVOicJOjj
rLJHgenitvG0+kvSMPQHICIV2T46qtGTbdQ0jkSaYhYnN0h1gsxr06kl3sSeyLy1ylKPcng3Zk96
BnEoiItffnaVmnvki4SFWVDs71CkgchJyb5b72fZSifnWlQ2vB0F7L91XrQaLHbyUmNPPbvKLpOd
dIB2N6UCL1IhgsSCcRfjn6eff0oXXjWf494ofQJTGbQv9jlIaukeUiuyDfl9UG3wysulfcvHbnZ4
8GguHeJpV5jgb/Rk2MeeoHOxNcb5ZwBcoJsYY+03bxxPF4kAScFpgx/AaLNygDF10H45wX8S98rB
ABrImDVT2GJPxse936egW3jMabnYcY3uyf/cYJ7A5B8vrPUgYpuvJcZk19/qqkUMsw9d9/MYaMO+
bkcTiESxAZCK5Du6b0uh0a4iSMknRO/gbmqT8V4cQ0du0PSk+m2kXJfJfT1LUP5mHmohhyMVimKe
BY3zGOc6KooesIODLaPSNl1o7S78mB/CmSDgKfE/qWqSAZlU/Lg3MRD3qeI1uK9c6dtJQDfmZlKT
ts1sVrc1eAIbG+iHTvZG/WNoiV1h9KHbMV5+NqEnoyCbs4XpTjn0s7tQSK9yHWn6x1SX771X6EOJ
uw69w/YscmIdAvQDmf4WI0S7949CofaUwfyGcAVM2EfL4cC5T6hZ2YJ62JZmS6UvmhsQzXaFCLB8
sX84p44Szhe41XtA7PiT7R1at+fv/MCN3o6Qnz+7xEH6/+pr13Pj1DrpMUZ4fCnI86ht0Y8c7oIk
W+rGjmKpGnBQLfSp12B8t0B1QKW6e9L4e4fp2zYVS6++cklHOIO+ntjFay0yy3cKyCmAWcaJVWMN
pFAYGge7qOfPn3k4nG9WqtZQT4nHG3rDBjgBC2wvRRhZkmbHv/jHeUQs7uEfkzbYN8yrwxNgxM9l
IlwrrZjpYJjIOVadcgQOv7OKW83DInGVHB6ungzlr7+IiNT53+s47Ih6WhjUQcnqPPOXSRwj8QHZ
rv5QXNzonyS6KWDPTMDpkeDWlo4mOomsZr0b6+ARFP0nTN9PGOpjBmu1VQiwkXnazM413ZfFajL3
K6M4mKH01wICXIkODZBASkThIe2d3cist9pPRpYlYFsbZAe62CorbAvhtpEC75GS125hGMMLmZhW
cfVh/cCTxOhexOLxf75s2QDXveC+MydnCcIgxjus0dGNA8HPIbcajedYDzv5G9K9mOo5+Hem0PrS
qppscXAcCfcgIaLHVCx4dUWO1ViaCp91alGXPlaskF3b0Z2fp2oDWRKfLPZMpLVygWpoJfesC9pr
lwZn0Byn9MXFX7KdkU/pqp3Ro9ArKC3ZCeuCGuKbAZz8rKXS9aRPmZpKcQ1MgDjko7nFs82kBCGq
RzjxMDjjUYe80omsYV6xnirxmGhTqJ36IJ4lZ41y82eODxm+03dSuVXhh6ffCzOTwUDnX9/jzF6q
CrMMkK7ukOL/uMz8YGWmiOXf4uJphTIRjxx+bq87EoWdOlNkz2kes/f40BYL5//VZFn75ospJRTr
IzJbx1SHecIJ0LMjW1tHXd0Rr0JBEjlvkMA9bI//gUkEY/4rQMlZR97lN7ppnkYi9r99jSssCAuN
axJHJ7Rp7pSeuW4NfzpjJaFYKbrZYqlgjCmVAR5XqlC5S3nzAcYp65hQdWIxIjZGkv95NNLUXRrH
3Pq8m8gSxgY9ST0cHP9SpgYxQEkpFPdulyBWPHaq6pqn2bRlH8uwNI+/TathBzhIiSbnjEgu+Xvm
ClMJKE2FiK0gNhkwTbl7da7B5ogifzhDc29gamWVcQeDohzxVFq4qGOhUJtwn0F6nN0mlscgIeOp
eTKba5u/D2w2qzImng0/SOGPKUeM5vq5eY9RFB/q3F/hSROFRGiC/YdBl7J0ayflBjNcJ2u0omH+
on78DtaX8TaaMdYMqdnCHQVWJnlBBuXQvR4g6/bMIt5XX0Tn1N32TqHoX3uhWoQbH3u++V3ThCSB
C69gU9tZRXpGFa7S/gDK6JlBNklHPqHwX5Gy7WYrkQ7U3CTA8Z0ir7zagD8eMarYzVt3cpAvBw4T
EkT75T2fH0K70QFsWfig+cFv3jx5yJp2r2s2smlWKV7euTX3IipL0uZhG39PbFaAP52ebH4ddxkh
Ym767XRzVi415SZsHDhLP87sl92mg+g7fmxvw4qRep5RZWu6vIsWD9QYmtmHlI14iV31aufpHb3O
+RaEMClXtVHoCLnxt+U4LGCeyG4QyPgGtTEznKjMwnJU34se7xp/aaUjzdwEtZD2IH+jIrv7gI2i
ieS1rGRkckA8AbXbXk5Ko1UJQnSyR8EM3E5rb9r9lb0Jvgtg6d6fDMN+R138YzQCrqzqDjl3DC35
Dk+C2f4KY1AACcwGw3TQjUV9FLXkoomoywLoIxmFijKaJTVeXPlSE2l74WRaITLOSMbqLzXaac3B
yFncEtwMBkC3ajW3JpeFmYDb2p6izwrE3cuGiqXeW/XsctTrJiF/65AffsjKQ2H/rRuidwCB+lx3
ibPjeH/IB01c/pw0GWYk+8oUccynNu92kB1KoNiHX414+ijLT8cr2CFvG8hiTvk7Z5oZnkeQB6Ry
HsPfTQpTshzjpcoAldjNCLGzPhddWb04oSWO2/UUvo/YJcu2P7Gj6TQKzDTNBhX3REWfDY/6pMAi
8bvIFAfmssCoJ2kP9ebZWNpjVDPaENGQEQipzLuC0Df97NlDUXh+q1ppmkNmmJZAXiSDuQHNrID5
t5/StChaZAmQlfNsLe2Jw97aLMggPfnkMAfIWWUVhOpFgdHfVZEtGmGjZYdQBB5eJG4Yb36t6UX6
Y6aWlkQdCV67F0JJ7Iae3GaQ6pAnMQuq5TE8fTHKwLcRw9iQ08o/ri/dlGIZNmD4VPVA1i8e+Spl
G1gE2bccxhwNTiu2GGrClmHQM+vKrHLwRT+VUiAmAy7/PM314IYobGlTU349yJ6IYJCWSwUw6wu4
ThRRic4DYp+TvIJjaBzlA+u6bg/5M9dB0qK9H4TUJB4q7Hf8BthXxN/OUsqJB670jgDGe6lK5Ra5
maWhzve2n5hEVN12X64Li6aPnGyMDF7YoGjKS6fOC2iniawbpM2+MeuPRS8uaCnJSrsFV3hx3x6y
kicW5OaNp0+WJ6EJ90WHO20JnShzO24o4G8aSFMPpVVY8vu0yPEHTJ/JAyILxHK+npQIWySHwKgn
KglYb3klL2mXLSJhGtysUBG5PvKgCLciPT4vN/QUVgMHGVU27iNwaTNRZSkQ+augOWsizbsyK3vF
ITOcPgw45T8/zsdkhvIMG4h4yqnnmXozcnApI+pgJQCTmO3+XcDrYW59R6wufg2skpwzUNsuOJLC
ELDfsWZU01Mlth2y3kjKs7LcCCvJGSiZCm93f8I1CtpkasJo9jdH1j/B5YsnjH1TSwt8aQD5qERu
MHCPstIl/b4FvZzDUW3wrI2LMqHT2VTGjLfchSd2PdBr/HtXaR9zCJV7asNYyU0sMl72cQ6zKYmL
/kzYeUl4OnaXPr/IYYTy3rCM68obE0Gs8QBbgZz4At/POib1outOmRR6ml8ppTyXhuRsRMcaQ6YB
nZcPw8ZXq+ueWS6rFdArxlJRubIHUMSjb4Lvop5gVeV/WPAMgG2qsIPUCDTgZhE0RptzowadYdwX
bajuxvfycprTJN64Smg2mwxCMJTTxeQXbZpmTaezomzJ2mSz+dYK9iwOiudB5r5kdt2+8BWlIztU
M0LJZhR/0oUTson+/bQWqks3RRL/lTwH/pwrqYPrW7kin3dVV+aOnLKgVi/pCKEeAFZQrg5/iRP+
SjmfhBmSgvi/DuP1oRV01XLYDG3m7HXjiO0bSyFWNmANQ0dV1O31PI8qrdpuahkDUZ5CFRfBO2aY
nR85/fanhoKkOoIMHJh3maVuBLnP0vjW337Jn66yhz7XMDMwUF/tu6jKtNXQBBwqOLQdpYWnxOh1
YPdzJ+ZNzsgHS3RjzHsx48nmT9x3bVNddFRd9BoSClTGsjTRyiyaw58RfCteQ/7k7nfL5gvt4GAc
Z2vIR1WdUDo5I8vrRjDJFS8+VNr0vHQFaYcHxHkIOg4UONt2IdvB6IdGP2WPf0tOC6LkkoXxSAaY
8qyjmiRnEYaZ5UlIli6dHHIH3X+5omWdARJ0DdeH0klXKtKr6AE3mNUU6UrUZgV1uf+v7MG0xnWL
2cswOzFqpbdBM13gMgkMSl1Z5Au+T3z9qUH9foZ0Eh+gCpH6IsxdrMZoPVC3C6O+czwfp/2nmpmR
5BjYyjqrSaIOG8Z35fwb0t5Bs2CZP+vcuoB+o8xvZ1WYAjlOcGwSwX3B3RQG6EAMpKUQs+gk6HNk
1S1Rsd7jrMLK/NCSCaifr+FXwpV/6NdqcZW66GBAivJEi2PBksRzl/Jlrta/AUuYpp9cP0BGFkVF
5X/Vqm1t1ayM7zW2y+WMUpHMaWmHlWbo8mAjeKZr0TRa9RulBbT/lKJ1DNmkQztu1FYW9n38/qSS
FHSuZqZvxoxe74c8z5riqbKC9DAqV1YPUDeSTnY3Oa8j+0VFygBLTDDkxjfb/wM54/XrgwgsIxuP
GnwLNOeC4n40/zacMmd6XI8tt4qbADzmKKiI0KZr4DJcW7QAuKXldmcvi1bSMBp2iPC14Fk9/0Qe
q3Vq7cJ/tUHzJEBjZ6aGGY3IN6TEaw6/d9T1RsD9Y/czL8wncPBuRvMrtjdkYY8Zjtbd8h1VYcat
5Yepi3mMd/WkyumLyBcR4n1tiAGEoe9PmlT7LkqKqZJ6DnlghL4GDYVioduQdcPlZpq6dsNo93Yz
P30x1kWSJ4nmmpkhFzPOWBDLbdeHcuwzKRtsYS4Bl2DFL+jA+yCDD2G7UM2eKLutBH4Sv7H7lscf
1RriDfVRsKgw1/CyGpDyTRoGuLPWvL/ujEsh7S53hOke8z4vyetpNMVMH1nIdlpU+RbucGQlw0WV
xCgCZK5uoE6wqrb/nBWVv4AYHMLCx6yS1mSFEh9jCF+T2QtYMTMGw+MQ8sI/7eRIyqz9CRsK1dBj
Y3AZHy41ZtdgB/UsCLii7RaPFX87qtR+Ep6SEneE8LDQkMFY1f2VyvDZBgpZqxJ0EBRQZLjqTO8r
Ae0YlOhDb7qIVRSz7hrlnmvglSvV6IN0/Nh2IRnu3LxXes2qEpOmUEomAor/hB74D0h/n/xvNxSg
1PL1ZjvYXM7ObF/re/Wwm0mF7xzZKp7hgObWAK+8wCEkadK22MIa2D/KP8MDq32etnaVNYu+sDEN
w7swaDwhgVbF8XJETV4HG2JiBOmlV6kbzn9f7PekauLV6hBx9W9gECo7fyoaBdLkrmd8jKHacmOY
Kv7ykcqGr+9nvtsDoMVnbRkBc5rfoNs+UN2IiF1iBRj0VGiqpLrgo5pUARBcBXOH5TiuQ2IIMSCx
XR+w5Nf2xxjfaiasJkY04jkbOF3RE9L+b/+EQcf0SbfngqnbxWuGc72O+Lertb5Fw/z2LG0l/BGm
xAUHq7Wjl581Q3Lsmb5SiAs9vMJdejAwpbzQnOhRJVY5RxrwLJlySKWP6NKVzHslKt3uHvRnAzJc
x/Xkah/4FAHHJPsN9YDHxxzkarjhRtBW/lR/XYa6ycHb8vHSdxU8jeQeYFv1CChn6pUP7QtgyGRH
RNygLjSIEmbqNAUxiwksHnw6HI3y9LJhurbDlLyqmFKhouhHqnpEemfQ6RKqhA2hyZByk/Y0F9WU
x/ni3iwFblex51C46/wp5Tq1AiEvajk75sWS7o7614VQT2nz33vZ07/CiPWf38OTqHZ9urgypMTF
RCzE0RTeYyeVXP8fZqJjYXNSpesmsJDOvm//hPRkafedbOWN5p8ZfC4Lf5FO7apCtMhcmWL9oSUV
bvxvPMlbN6CeoIoRi4vz1VISTC2VwHmiiu7OXQqZzJGQyGTOnihgb33AMVGuoy36xjUhe08PzK2I
MX/97q74C+DOsVkqVRoGwE55DbOQZPIEcziSe0v7EAyLOXh/13wL+pSvFCgzQKPF2tKs0n4/qCvx
U083oXtxrn8TctM5A634pXFTxAWQOfXrSWflDz3Ty0mvV4j3tA5GeSgOwYM0isbEa/ZAtFE/NSSF
xXylCyQRfSGGqiHfw7pMt9mj2stWRliFp4PatVywAANVPjXQkYKo2rxvfKZ7dE+IUipvVcE7iEkY
WLAs92CAyRl4Hn6px6/pyuDgpxKS1PaIfOexwt5T2ruRSn4mwuiDp2JzWMtowvLayhvw5dozIErV
TIMmr7Ywm7qp8rjm/HjBkwSbY4oQZIexFwCWT7cBeeP6qj/Vpi+rQXFgyGAzCEFXn4W8XmP72bLz
MS65xOAZcCcViqGzBGxFF9gIvB51yxFZClvn6rqvzpOwv3+lP5bDWcl5RkHf2VvcZuxd8XDOq1Lz
MVMcnz26xkPup+vdFbG8PPUSPYfJ4SJbFJ0lxH9rjfZkZS71ZTbg1kjQEHwO6+F+3r4bNyK98XpD
ZgITArtGpmRmzwWCfaJsJyDJNLUD6BfLMVSAC+DTpHeD9xWefHQ+lNQRb+B1KtxDJgoZz42tQ99X
GRhgb9ztBRuOQDHKplyOuLbU7Rj0L49Ri2U0yd5YOakU91+WLUup3Ej6k79KcxtpIDb4dTFd3O2P
cMPWSGTrEqQ7lQHC9e5HZsKM2w4VT9MyFUwCEifLZlPuAQzrwpw16D2AtSznwWMG4HK2BHw4snxq
0S9LlpDJkHYjN8nk5L5PW9LJoI1lllnbesOWcz+va0U5RjlhhVrNh9UZ0yvBruYOSeA6T/e12vV7
fXrv4R2sG2SRWdk//oXCD3dnaFqoCYzAs5Q3wqmlBSCrmh+9H02EALh13AmvSEhcxTv9CU28Pvss
dYaV9AYfeMGEdLsf0VinQt2cEfSDfe1sgxG2EX7rXF15HfJzJEnH/SDh2D9BtpvZxFFydBt9U7gn
ab5m9sm29XYrzMPP652j+tGY066EgwcjBJW16w/di/o8a+/zbjuvjSt7Uy29+B87pLdcccKiWmK/
u/kboXs5qPV4LMcKubugCZecd0Mpy/m6tV6yOS7mkoAFI1MkHmXLT1QE2rbyomK7LozUYwk1Z5CU
RenaeDbjGzl5saGnfihS6KZUet5TCNiXBL9Bc9iFHde7Zm/jRjHkpf/t2SCVNbTpZVXouT/jGLcI
Fo/RGGPjkJ0xHb5Rf0FKhStvv0unxTuztT7Yc7a9gmmJvBk6G0fLUtapVXCc8RoITOuzAo3pMZ8s
ELjus7rUjNfmIICKuXJuFsO2IJhOZ7VDEBshvPgp7p/BAcc0Cs3cEhludjcivqt7ZuapT2g9yI/L
DZxVXem7TzdSNhYTC+CY4/+b5zqzBF/uTyHvvUjnaMeEZzDZcn794uCyegfKTRUWvxTw1qZGrRC2
IWETPHIY2midVLcgwyVYB+NKM/x4m+fIEzUvrloZsFkicAunk8IOEMchdk0qzzgjCyBfiOgcQ1zz
QJT7st/j+TnMbK9hNx/b4Cmz2GuMnS7pNnIJsA8iGdGEtsyHOtn6YzNCpm/X7eg0593ty5QktMP1
nuSKi/Vxuj/1jHdmdS2A/nDJ9P2eCHeAVgzrsDfFyBl4cfIATTZdjBlF8Ex7TYi4ZEpbsNuGtFXL
IQ4VQDqQeFoklTmYsBff5+6Vs6uSCm/ev976rTKzSZUzdZPdGyurI4Zitm7u3/AG/eovve+Tlozc
2jJ0wvuYq2q7H0Y4+KZp0cqAYRzoHrToTPYpm58ViKZG+0B4OzvroxvtHw23gBA6ccyKzgDiVy/1
vnELE7Ylf8s/F3VI4HHdzpXWCo4QMQQ9SKysVJsFuzzg5hYfHxnt2jYWZA2lHwZFK0Dh+gACb2Ec
ySnyXQKU6VmHfHuRttwXfuEk1z1N+6fVpbc+M3lNvQ99iHNGyW6ljMJsOdxXQj8Of7B7kk39zS+0
pooGydz9T0a8sC8rWAeNrhkCjpj219mFmI+SO4v3sm7w9/xHV4RLuHnBDVesLcGnKFwL+Zo2uoMo
9wClZIAGLyryveWbjstdM7115ySclBlJ72GNisnK6SFTw9JJ9qT3CthSZOqu6vkgwxANKzewvAPT
hz/qjzunj0FxKZ0iEA5MGAYuIUJBHC8qY2n26zCk96VO2tqDIg++a55a/yF8Op8sPW7xERdX9MwJ
t++Pd7hNaYeSA/aRee4oGOV58E+5F57F0aVu9AuZNOhj22/BJkCTTB7JtVr9kkW/pGafB11/9HkW
IhcbprMc9wzc+DN5d8OP2Ku/w0+DNpi2WDRQZkmCSDzW9jTJ6PrIq0RxtwBz3JHJAPSIJh12b2iJ
EdhuTbuqWCs8ty2kCouCxs8dLY58ogEBk0tOw6T4a/qq1qt+mRODuCxDmHniV1gjJzCdbRU8Byim
9SQSNioFBgfUVe9TqSmK6xw/qF+APuZrobGKkzEXD7o8C0eRm8MW4sC4hqvvAcCkDvtpKxY2yYEz
rPfY7HQVseIJsxDYimLCieQFIiyN6m/sq2yY0HujevQ4/YLBpkGoeVYDWv4XgoTRUxlYqs2YJWiK
8k5yksn7a7dB1dCFhPbCUVa3bK7PNNrcmC3AWtFftM6u0keh7KxXS4U5TZkENxr/j30+zRqsyS3O
iOY4ZlheecWj3Mw7D0GVNGENeNoWjMRyw5zfITTX1risqaJaXIvGcwqCHc8JKADe4UWuLQFbGHUQ
VTZXAu84SlOomXjSu/67EKf+EM5dz722pesZnjhAU6pMD4kmMPQJ2z9LTs4e3Yv/zCxXl5XfznyB
/FuvI/HZkOk3J3KRRTBLikibLBx7DttpQLe+sf6dKDH+7uvc1F0ztHHdegNd7IUk9a/Y0g8sjiF4
vEpobAH0GR2pwJvFlZYSpki9E4CVS+CQPTdpkV7xt00NUxbJ3cpC0vYgbdNm2rccXM5ZTsot+jHf
YEFw7ULKs0x/0l6Q3kYr8ZSvqZ7BY2rg3euVkN2XVRQsAhO6dzztpC0AwGikUZfSmPtgomYOYP0q
kwmLUMu5v1ZVXXxBjel3y3EZznOuet3VAHe+vCBXO+IiBIrYjuEY8sw6Z4yg5K5S99zySxHWxibF
iC4/cRpfwM38KPzCL7uQrrOPaljkudpb/eijhw0krZ59G+G9O3ou4JWIt8xEX+ZUDE8RPopSmQOg
tVyGfidcgJeGHJPP+MlT7MX9ZIkmRetPxA1Fs0F2YNubnTXLG/lwkhsxxFA6/su2ywSnoqV7vYOE
x4mbKassk+wRBXG/MErzrw1a4kjSqxWLTd2GanaCoJpAVQbAvJHwR+mz0B6Yr1OK6HwpRMw/oARB
Aj5PSJQAlmXuIhl40klUpRjuX/1g62WcN+a0moFCX3WFwGbZWEiiFAGCP7Ug1ZPyKN7z5eEdUBaP
X6F99aoZUrmFxkLiWn7EhNhz5oL3IFChRt6I+g7E9k+9fTHdBlb358INWQh9R65OtrXFskqs/ig6
N8DJ5OVGdtaadmapaiXSDIZGFdqnK1ta3zTmDtvKmigbCddG4vvSrXt2bBohIVvzF9UNoJVF4MKL
d+hEdLaBozet/HqtUW++O988mYtQBkUR3SQmWZQ4IDAnFcf8eU10O0UKZsWw1vWaPtS56eqZO5hF
LPHmdt0Bz/JQpW5/yUy2gz/EDvH0QgK+azPkNNW1OTmeVMnM0OiVUNlGW3XKreqVOx+PYQDdF076
GRBi6klyPIRRB3zL8dNReyEz8MDoS+o+vUr7kgSLm0QksPcoq1kT1b/fFu6u2acoOk4n9Ww9uHMY
snFPYLPzoolEIklLgLyCpGkHeAg8lsSMV/nuI2qiZYJPHMfTuUfnpQgLbdj07raGSyTgdS4h28mb
lq5AxGEVs6L5iujkuuxN2ERyb+tFY8Pc2Yqz4m/yp3Ingae24otdy6yXS2+H9RW5HHIN+z+t0J6i
cZQaUqFh5mEMI2YLNPAbOJ5y1dCc1EA0zy08XWB+oufkTo2Gl8NVh7pOaEvIYVTd6M5NlfFDkHuf
JoU7DBprMGxog++fF69d0zf56FXEeIfKzF/9vbBPN9yQj0l7XU0QngXz7HBeS4eTHWNn310k/h95
j8mfg9ih96tA/3+DptAnMPlEhOkP1CiIPYLAt8g53th9xabbLDHLKZ5fW88miXyOYVXrfK3Tl4BY
EJKeDHPcjIbXU55hewKCdfI269+rKPDJ5yCbAoOIoeIttevGCZ8cWoaKMQJzWByBh+qTZFkdsv7a
FwgRlp6ezSYdaVjy+1sCeT6dM8dL91OewqLcL+e/erD0Yxr6MgrwSgbWLPRA9YgBE0kAJm4tcxra
fWN/qszjXP2kkeRVMXq45dZN7g60xSFOH/IqdnAFCwx3Vx+fj9LL1dWT308+QbTKvyax2ACDLlJP
52D+xjXMjd9UoYL3YNYkl8sJL/73RIsvgmnBv4vKwURgn7m72lqZUGXIkkCoj0xEyL94H5CU56P9
scK5uEznw6JfxnQTsyJ88hGw4O3Res++hYdqR8uvxIMFYjoPRUcr9jzBadKARW1pQPDGNM7IZYVw
JrgDJ7gYMHiqKWOOoaodRHMqY46QUwvH3wfGL5BSUun9nNOTpmAhOxabotfYHPGNRaCEOUQXXfUV
Xcj9t8lclldyS1AOEeQeD03XjQ3SPiQxfAyFqZd/dgZrnJdkXy8ILlML64nhQnHaQQ9V0gO8WlnJ
Ol/NJrBjzQDZtjUuxtmZWkTPJsZeu/eQbp2LCNmgO9rxEapc3xZsZ7axqdNSSzkwL4SqnlT80ulR
geNTH4qDRh2RqOVjjpqh16tCiNif/+SKUIUPTexh0J/Eak6LjvJ7sp7b9oCzzM2kH4nI0bk6XlC4
ewrVhxtLSuyviJ5fSOmk27WYuUsDiGPoqYDFu41rUuHbnUlpuWN05FBGrRCY0DM2sQCheMl+ePCx
OgKINRyy9EWNs0qeLeM9qqamusoaFVFWJQuOh0GbnpsENgQl6FphKNkgkv0b5Gs+bHARN9EhqIaC
prZ5zCNj6FzRBsGpVmorzfOgh4BeGrY8O7/S2CSR6q7ebqk7LHsKNwuOH9AOPzT9gqTskXvXGvhS
1YmKX9YbUd7nlQA+I6GrKCqUIQ+i2jN5EGlkwPCcFPdJfAKXIq+9Y1/3tmwgSUrssTw+Ct31FC8H
Uv1nvLGFc2WW1emozo8FOEZBemf4AV6aSWQ1DLouANHyl9Qm/EArFOaGRs2NP6IWmFJ1xtFb7dwb
kkYzzzXrNbu4yE0vUuvvA82ZnjDClZ+P/f5XA+HLJ5eHtYOpcqdi/qafWAeAoG5jqodKS4cmf9rp
v4CfO5x92I/JJe/Mg3qbtm9vuGfUBrNt6TuVdg5E/un0OaGrFGGZFy94GGCJVtmXWMeDNQpr5TmD
wp/wqboJdUkDO4itP0HgXlRiP8HeDatJVjR9meBOXQDyz9wvuLKXd419WGFMBLoiz+evgbK7GOh2
UNUvL7RO6SVNqUR9OgE34bWv3HXOkIrsq6984XYMWsVP+mW1u8KRzZp/uDldj6WqliyIoRJZodw7
a/+nb7CPq/kYAZt8KLEy8G34qOW6bNZNB26ekgLT+3DH8uL7/XR7e+Cmbb66bbj1cmjXeIKhNaEc
5TX6ZIvqOjs4Shc48P4e1962fHO7YWdD1A95AreGrfwVgdhl8wdCDYzAgK89wSKo4r490YYZ10nr
70qT8i6ZR+il2NMpdVq2Q98Aw+grbLSgxipW522gPi8Z3putJqLgQyjIkZcKur327IqfRPk/0X/r
hNV0SCOFwPTOqywwPhMSPPLY+WYBCIrhZ7mM9zFrDUgikbNwmXj8uV2RlxoQY/T1dWo2efaqGyjO
wqhX3lGwy3CF68tAQnJxFHsVd6m2IImgTr6KbS1e+HOzijBjKX3vCYxgt3IWeP+L+kjtt474fMGk
81ygnniaEUKTtVhuyd++jewbHf4gjUdVE/f6ls5tRZi3H9Iabs4xIOdMFq26ZAXBTYNE1ASKfvTT
2IhZuvrFF16I2OM0BIAFhYN0eeT3CAh7V3EVBlOD82vGTzDU0O9ITkHXd0FpSYJVVFceCkuapeWz
O2inYmISmdMtkUJTF4a6LovEdmfeXaX8EMc/HidMMZkQi4lTa5HyzmAra98ksnxowt84Rzpof3Eg
ifvRhf9Sdv3xxBJ+bAN3jGsqp5nPHRR1SV5KrBLg43VxLGjwE/VXT4xCHIipPwsx5l9N0cWXPXtg
Scbkn9QRUCaudMJThRX37I1QTnkVdpsImDcWiEnfm2FCJPjaqW9E54il6C24e/ZG5DpjdyTyysdL
XqkWz0Cwwoa2nIAnA0wlI6TZMaJAPOEQNLTiHdn3ZjHbzCmmJWe5hzuCRlbAs8LfaSkp2vRJn6HS
HZOT4w5uof6jtlRKCvzU6dupnpFtCA2kEquswrbJI8Vkc4FgdnazOi04FeEYlP7+h/mhZtUH5Qf0
T5T1NHtIibvuzfvmqhHMHVjQ4UfMiibYSvxxqsevyDv4rk+0lOpu8a3hg9YvVViUY99qhYEBj2aA
1rJRawaKQfGf55VXVq9Ry5kNeQDDXmKgaVD1RmETYZNbDhGbahc9Tu4xvWx+fEw6xoIOgpbwsSIz
ggP3gcCEPw/wuI5s/i4K1scdBCHNL52u/88eNrs6cOGEkbnjwJT0zVoCQdd7jz1MHTK2+Dgi8yQN
2v1T+DK/7i5qf840iLESnU7W58ahOCbfCvWegtD+ynooYm+qLF80AtnWk6kS5i/4Tvernwe16TxM
OItsmLymBPW/SxRJV1XbCtWSahS8UWLI9VEXh8aMWiPghF/UKQf84hcITmlkmzBMgsnLognYOWFA
L7W2qvqLRBRj20Y5E6QPmgDq283HEfp8TIHNvw8UtlAdt7TEI9KC23U3BGi8l6GNREbZtFJCeAVd
fsYUghr6XvwttFdtyb8/eGHXXO0JQakisLfO7k5bs3EwhMXRlqO3/FKBq59xGrvBbS64PNeqrovO
wqxApyDltafbn0K0GFd4w3BpccE5DX0tTeKyOtjyOqgLWp6xUfKn08mN8d8ql1+BED+mljF3bSfd
yKKATHko3iOicaskcyM4KnKFtKJVqQ6i7DRe+LQqUxtbLC+TnnAgWMDTOh9+o3/JeJcW66IZX7ve
KexCOKwST/3YIsgcflLh6kKHApU5uSMNx0gJpk1e0En/ns66L2IPeA9NQoajqCAQnhaxGhpqLLAn
xulGWo81AOKGrsn0FDXsSB64cqgdYZQlKBDFOFUSHI3IdrKGVElSS4PIBAP7q69C7KHYqTxeiOFP
K6BH4jOQgDdhyt2mwdHDrQp3LKkjdcxrRIGALKthKoQWSv8WUFakJDPc4Blf8jtJkLQ86GKaFByt
wh97mWPNd5zFR/EH+pc8wNm3L5ePLs+MlaZfOxiUlgpw5jG3lvKdCrWBK4aO2Maevky/MwHc1sfs
j82OsXabJcV1RzBNq9/QOka7OqAomHfit1J1BBO5dwNcXkkUQ05CIVmn3U5yUsbm2aQ3EvZUUPwX
s+GwJu2qybNbZzxpI92r0/IgLKVqaPkmkK5Cxivq6Af4wLSNVGs5JU0jS4VWIeBQsccejKT/vTsb
TOuixG0QH6lrUpyOn6+xtuyMOAKlxNwgU6eHcOshQ338/60SgZEhjKQpSgfWxvkQI6E/7GY+iMaA
ItexXNErGIGaBi6F+KjLxNTX0FFxpUoGpJVGw80Pm+rzJmKqpLnOzkJ3hBtNhs/+mEQwBUZa4fo2
sKL3CdiG4ktevRWM3HV9hjFeZryoF4xck7ikFMVaVUckTAsdRh4eMlMWV+vc5HrUrat1dJJczkhA
Uy0B2WayAtmJBufx2hE6S0f24QvzkElxpBP/ng1KF3XchStOUtTskxQxxVc+MU099Z0dnazSBhHN
IaQk28+8xP4fyYfi5Pj0bAfBR/CrueMknEltZus+DY0Uaj866+tgWHuHIbmKmuqJ9B4/ikrwT4Oo
YNJ0AZqW2x5/kPxt8Ss08GTRAqjFT7L/iaP/tbjkNJzKLPxQLnxBJ8uec+7yDXplHcafuRcBgm0n
wgxUxwHwQ5Q2+27YwadJiqfAuiG+uwTvtqvZBlDz4Lm5A3O/DX7bVW0tjN7q3IbhH+5lARPEv5JL
uCkRBnLcrUHO02uvYj+d6xMYhN43FDZsGjqn8Iwiw/adBByZBLxOrUDdAPoCOTM4hCIExEoRRBPs
IYRvgRJtdF5kM3ShRCW+sLBd2d50fvF3jMPI6KHH6K9Bbt5TOoQOnKfL7jcmtZ3mKqbeijjeMil3
1mUXfGrSfcv9MUBCQfgg2URB12um+pxySICQzm9d6/XNCXDvTLJV2yh9Ku6kACnKuau3vSgtSROe
mU+4qHj8oap2CHABNJgheR9GBi0fb0VqMUvr4m9o2IACLXpI7oDz0GiQ3HqyjS87ntXH6vZ4OUZO
J+0F+EBviPl9Vs4sJMLhE0NfokvBOSDGsTG1S+2mYPdo8lmKdfOTPQr71tMjUfc1Y20+kzwEPZRU
5hMoglAlF15JWZzbVfQIKMDD3LseRHxFFr+xZX8aer/v+Bh3Iqu0HqY2fdvKATc86hLv1Yoet7eu
Eh9hbkHnXpGrzVCkubpPqcJRQGemEA+3xwvaqoL6isSBOc5cOIRr1RIUDUtw6Vb7GmOn0bDRUIaH
P5YUn3RtuPn58ZokncRt0pQiLlPfAuiPPPjKvCofu/Wa515FZ/arIPK2gXO9SIyXg6RNzoHqmEry
LQNhxruFvV1fYnfCRru33u6i1zZh/2jZaz2DFxNpFjzTWIAVYzWO0u8ki+CvLwE9JBFpYUzTcWW2
D2Rfb64IAi71Sz24oy1hp9kqCSL1P0AFVMMyvC4RgkLs/qEX6WslZEmHC6N6vxV4WAevVSoZn44I
w4fCWItjgWPqn6TNyKiZBpeiKMNuZA/ypNsr5HwGvwf9UK5lyqT5YTF26gzci2xJaD1LRzNx0ZI1
0QQy6PTB4y2RY2tbgvbJoF3Rh7eHYJFgbuftUP/FoVXrc/U+BGnfm5nkXuqcSbMmouEIuEks8zIf
L75VCoawRUA9XpfXJ8biYUoXTi8lyPPdJZ8c4Se27N4fyO12kCBLcykBSyihVVn/nVaY4FdaF/DD
5Sqdoj9RlgelVPPpHZfDCvyT92G3hHXswWQ1zHoLvTLfvL3rgMh8s+0HYacAWHSsE1slbI4i+hlB
IPO7dLPu16fIs6LSnJrgY700F656xWA2f+hnXxdPQ6/r2L12+WZhw9yxy2Q10MR/MNXM8K+h7Xiv
5NBjC2VPSuCBz0BX7G65V0KQtSWp9VfPLYP4RWrm0CwSwkSLFeI2UZnUTMk+FKochqX0keQ6KFuj
54WxQP4n6x1E4qBlRGaOLCLbv+siGZDp+el1mC5xdkO107N1VapnoQ4z3WqnEcSVBu4AZYheWtEr
4wndr4CB6dztP/AY+MmV/BXKxh7Wp0RNwXF9Bg6NjtyestEUMZv/KASwnbMi2peLm2ky32q3nv4F
1GI6lf0G9cx2o5DsLjx0QvGr6Kjmjb+LBUAh7pYXbizJsMm7UJflMfnSFxv56Kftb8/ouRHiazrR
HDhCbrrDWW1ppceFHoghSJ+mnwU06km2I4mz09h0ZI6wfJXzNGOpUfW3XeRXSaI3nGXe2QxEwT+N
InV5MRFK+O2mXau7kCBXciPqcQ3kTR1tI8RkC09nJbtpgqSKhhSDdXu+/7Jcw0plyojUpRvud5f8
3szgZVjfMHF1L7cgrHHSDindQWo5wLgrjxxx9tLcUmQoWy0CZkUi44Qo/lqWm9Q5eIUuHm40Y2hK
DZVUMWB6GCn6vQpCJGg5tH0dHRWr6V2eNfLyRBd2itklLUh70SNe6T+Exak3qwaGVUXjF8ORsfEo
DXHnergr+RsWGSgD7JRtWiq12K0NIDNUliSXMO7tusmR6WH/hBB/P5j/Z/LuWhJTPHAHSWJ954S/
4vQbRUVYRv11x1NPWex5HX5OPCImHGGToQDZEqKeQkZrhW9vskZVDOycOqr2nRjWgor/almHFGE7
oScHe93kjCu2eEqPgwuBTh6ej353KMD3aar0pK3cGR2iaDuUgqE2vwLi1vW8EHo4YHR1WHlLHUof
M8nmbGFIIN2KP36vR+npStiLjcZImRYoobJFGSqzBXDIKjbpHNRQxfxHMMVj+kvdJB8GTXBdj1Se
fcYLfY0IaRGj2oOs1OPmqwHobgY1XDzKa5zSFtfVUXBB4ogktOakyQztJFOTuyo6DU0IdvTBcdyO
S3xDpzhixeiI2pQ09wizkxCoUqvmPIWixljr/Gvotz8v7vl7R533BsSgPdj4nSdFZDKeMgEbkghz
SvouKVkXsdEF74NEUDaMNWOb7R6KoyNR9jj0b7d3SI1BsSqUvYBvUAuUwv44Pm8Vf8//onYMk9VV
IBKAfLKEoJBRDZ6GqAvJ+UFDJnXDZs9kYAKqih+clG0yjbhD4fJ4A4k1VL35o0J6XXDZqfIZanV8
vM+KDAj8yn6GJtHqF+elq3GKMH4iP+uYQ7ZKdPesumnst/GUjce8I6zqs1p1Ze/urix+GlIX+wcL
T8Y3qcIrqf1ydNBV0N8BKIy2wyVRt8kTWJ76J9f21919qFRA2zvGo/E6/SAghqDEIVjv7s7oUh9V
F2E+ivQx68X+/CLRhVAdcWCMqrhiHQhaclxwKS3oZC6ee4GZWX6G3oS5ghw3gMROeiYkbP4P39zX
qRTLamRLw/JsGa3foSdbN7W6wNKayyEI8Sp3l3KmCVmcu5qtzpxSrbbebT0hBOyUcT5nCVX79vFY
mT30SHMrlglCqiBHcsi1ngxJ38EhlAgjMNvmTXL6v84MOwOTEah7Dpd9vGj5FaODrOmZxVVMe9y2
4jd4il8h9qxNJsP95ITDaQ8PfErki5TYp8fbzXnijf82YNPhBP3EZH2dGTKD+KZ4dbRQGF12xbcY
3cHP4/Nn2/D5hTM4N69rFTqwcl4ZuITJvaTVgn1DoLbSGoKCSuv8oWWR87wtsOWcqo9faFf6IRF8
0xMS2eDiDgUKQJImNWAoY7XHOmQjpLyf+5BDL+J4FGMZX8fMxHgV/S5w4mPxp4wdq9WjOL7HUIud
GBgMW/syTCKONZY+eoBK51G3POZZArfqlNXr8YcLkERm9XBqhBBd0AzZBt/Ut0otXvybYDp4QkHl
lnSzPQxH/FCLHljZIv3WQE9Rz30Y5orcOoMqu59WtCGJIB6R9XcAS4TJowCUnOddHXgDKNM02dQG
NJO9Z9O8rHk0GCB3uOI7e5mCj71ZJYpRowNUV/KO1J19k/Xhi62ehFzORo8u9T0clcJ+ZGLt+RaM
rinGeEgwyqvBuReEk5Ac8THWz4TazzvXPbz2I1fPo0qAh9m3kYJAGkixgAXNIaA4WMA93jaICx8Q
5Yz01G3KtNbjM5NeRmSMZ2frFKavHA9rBHKtl3QIbH4noLyt2F1VDOK+n0kr0FVezY9uKGyQXZEs
up0drtzZCWEx4ARymiPusvjilK3XFXbSkm4roanDnw6wv++JWUj8OTBzcY256NbTsIgYyJR1fjIs
Q8cio4/5GVelxYgVNaHr6ECm8CWVa23wY4SBzecYL2BAJiYJzl2vmEC6kDd4xrVBZue1dinTSPDn
V5OUHHhJQ7TV1U6OHj8xgHmkZwrxU4s5R29kljJ0uNKf2OPxtN4la6gagWnSJxJgxO8tVsWrzkFB
9Rry7OVp5o60EmGWaBIa4aNkhInGIsV7irkCyM1x/PsoEcsSY20a6z9mzTOYnXont/TvUTCqnJbY
FzAaLnXpsKvaqKhRMQg6z6xkh5bqbPYDUfCzBniXRpn9AnnN3nz2Nn7OGLgOmsrsm3Mpxt7ykCio
N6ncWSLY9qC2aA7Uud7hpkqkJeV56u+GrixNpRPZjf+MWnme9Jx2uyNxVqkIz6nPJGKN/j/OnawS
JlZMgcZayCJW4/TqUicDzzS06f+zs1TI/Kp1/zc5kAQKQrCHKna9oT4oXTqobEACS8ht+UONvYmK
XxDmXH6cs4EqFDQAlhVp4+lD/I/AC5PC2hdC6nTUMx+D9kRM/i7WokrJ9ouYfaWzgO8Ij7IDs+Zh
S6/if4xr1cuYI4bt7VkZJWkPmcaqvK6Kt9NIQreGicpDuw3xwqZEgiZfQYsbh3dVDEFq1UNiRJVi
rspyuYXap9giBYYzaLXR7xDj57eUxqaGvzetP0M1nSuNUxZA6zgIDWeWqY3xqU7D9X2XnorcbGuA
iqo239nErqkmod97AeEkVRkdIMC+hbkiHsc76nOlP6uByKztByf+3CygLRbQqzxV8iicgzhxvEMT
Z6B8WjhmMx8qDRbKUgguTaxGlg8JEGTbUjLATdqS7DBn5wZoIPDmEYuGVBZddaCvh7sW8SbW8GfZ
VPOptSDgiWqkOneaQ22BkSzmu3cMJ58zsYB7wETtWVMqM74u+Q5Wl4kIX9jcXBdrrljKngnKPYz+
PR3FsXN++wTglGCpzt5QAxnFSPwHiFTnxhOT1M5YOtlm4BGfIk0/bUXPj5lMZ3i/BPvCC2+ky8WR
0M6+/dHUMB2wgDKmNwF35Qe5quRW8QQRGCrgIPNlfDh0IK5aS7/xWxFrsJu7eZjBjNzk8iyNRDot
kWfEG4xiTW6pstjZZNW9iAykclD9MSCWotTQZnctrY2kLs4lTqmSevPh0gDieICSHONcCu1iYonU
c6FcerLTLKSylxiqazyl+fvrdoBu+DLMHVm/IKvAJ9YP/D8Bt9KrXzKmUmRZglxl6k4LNEEFfYPo
BIsYysGK0MfaRbEcn7rGEEq8hGmJ2q01rK4CbAuGQC2IzpXIW2A/E5D5LxSdrfNnXXVF+teLRbmb
GpODwPi9oR+RxVwk0w7xs9DlSs26rcSA+crr+xpDPKJ7L8MwgZsbIk29fbq9vGq2E4jHTVXteTUM
j1QZuYtlucG0gNViX1ePptU9pzVXrIod4rkXeRkMFWIRYYkI4KeLBHr/FNvclmUvDKD8HKWEoAKB
s7P7EILg8KlctyTGAO89zy8J67/OV9imq7a9z3mjTbYsak9ijoAbeva9d9BMfCxmD1NDFu/ZgDfD
CgSjUY5ehJWGXmGPDbj2aDQLsaBYOkowNU7Z/cOUDdHS0NpO/EQfB2Ln0mx2t1DAVQccUnKMdwrF
u091qOBOGk4z3JFM6McBSF7ZeYAJgs9WnRNX4FldJSCy58wuIuTRnjMq3GSG1KGAvDAjpOF5ZeIE
fuCBzkYjt50kr/hf6GrPV6+lcxDcz3DU5KvoAUpPaKFULEm05cuLgk3jBqHIxtVbedJ60oe7QVrU
v+D/qWtrH4JeN9xsHggYkS2n29r/3hQgGJZD2lRKeinBFKc0HbcGKSgWb2tmxyJUbFhAJSgebDOw
1C1nk/PD6vu+hk6uXuC38Gh+pc+jYnh0NczzW36RIM+wdn8nipGfCH4abrsg6Snlvs3SCS5U9y5h
8ZmyV7cQqYcj2HiyQfREHHTZ7hAPHlXv4J3pegwV3IYeg0ct5BKJSGKGI+DsEqqhaLHydVyhEQpH
dqIGYUAV1WjgFJXgwsYGah5VXuftj1Xqhz7D++QZYlcMzxLMbqYE9c5dariwkE62VEI7kxcxURHL
cWZT4FTjk7ul0NyC/NYym6dlwceRO63747FeCHj0R2h1vpk/Nijg1JD0aDt5rgCgO+5dA/j0byAq
5KhGPP47EH8DPeN+aT4vpgqh8ra1WKGU0TzzsAOLmZ2aFJdye/YPZYhLMCPkTXqFjv45ijZM+A2h
Ni6v+HBnPEb9W2SHrsh423ouCiouwSb5dGQnxhSQE4zzMognlVGbXXCr2mwuQ5GBpjWTmFNeK4+2
7AWC2OarrVoYXn10wSWQ25EBrrXdRkXJfN0d3Wbv2MKcUSHEiz9W+zQn6CUTsfACpxvR4yseM/O4
BaFycQbTC7iUZBDUzyNyLEdL7pJhmog7nUS0jfwGKdKAaG0u/azJt8bo4Hs1XmO7pxotmDpytZBi
qYby1M0Ces3vmnxj0UpgMHJbtOxC7MjjZkuzowa0lycu4auikhL6+iLP2wmDJgnE2TMF8QUqxgky
61jirzmhrzsnMgAnxys/FURfByHQzp4mGYLa1RSfjeRRLC2cMfuROC1bbCfgPh9fLziWPABTOZxn
/IezhBF1zhEl8Lqz4vRzOJUsNnWuMboDctO0gxqsLxtxNR+E9/YNTjQc3MXX8kDE+1CAlAjxX8ym
hCCfzOFGLSQF35cW8jLXajVq7Wx2h3ymnfMhjAQuaDowl9gSoO87d4eW8u9vv+2xHMurk/kaz+wj
VWCQan/Annkxo8zzjpglllSWsHL+zzGDwntgA6Ee/Qt2BTewNaEdm70NgIYVQvp+Jw9NCtYXEBO3
18Fs/lKmpQPdhlU2m5ofmHJPPbeClS9CUaeuqLLU+arLr4/6P6ilijRvFuJxhu7gYPDlwjHLXJTY
yIMabxcZkWa6VB5E9uGK97GOUbsTtTbeEsRkGceOpdQHQfPASfXWR/b2BXbLqt9f8COsKdXOGIgn
/THHLbFWhnJd6vlE48m2/+HhXr7kHZ26MeiMXO2ioctfo4DIpcDnVZzJsp2Lx46PAUEjN1uByLY1
0Dl3o0qtqXzDab8jn+w7SXsqvv2n+F/CmV2nhI3mFnvXrnmgBzjPZ02KvcHVXz6bE/mq+ZFoxXRX
l+L87XsM6cboP4cQ7Lmoi7L9hPMGSaVkuqSn3+t0R36IXAsUrRxyARX6Rq1lkpr0SFV9g+MuTW+h
WZHX6iChnCKaZF84ACFNcnhuEdl7hzwgmEV+uiGK4TErARg/m2J/TEyq8ehKLBa+ZNTkpAKANsOa
NCompKVXEsYZN8seWDWoc/CSFP1WtH8dO9/uwjyq/x99ZD3MUu6ejOskFNxRLB18hxqflYMBW3i1
rqp+ZHcigBmtvWqH1FARXzbUxQf6702WO/T1R42OpreIPn1PEhK92qTl6Y0NEQGLQIq1IBt8sgk4
rNgU2WzgSVx4EIkl/wOzSaKlmpLI/Kz2cstb2JEgQiizU+tg84aLh4n089n2e53Vd4G2CMJg7wCt
8DmQharKqB7EiPGqISEGOOfOu7m0UtmbQ8wWtSKajts6c9OfdVsPEjA34i3etAUFhCf2rqX+rfQ8
qcuEUDxdkVJGyoSzC8E3m5+BWXWEpN7Uhv0OtAdlmQeq2iayQ0m1XoGXY77jAyWiWiBhRqoppGPQ
mLb+86KKIjqxLUbtff0TM+2IXnX4VuEIOzTIpmx6UlkvvstjV7EzePsde3FCIfW4A/NKejGtZJtT
+yWavFYP/obbu685UcwufRGVUb2kmkx7qTMjEleLcYBcu8X0ILTfV7HX8u+JFbJ/tMyybuC4n3vz
dKRdEg+EEYzuUT3xE8NEGfeZv5HJUlHdmazLEja601sx/t+zTpj5/B7snngjuSKQkgFAxC8MBVHf
PV2rSRdHu7/Q7TdbZUAtGFmkpqw1FHWKjNc4apZW9Ugi4URzRLIPcADbR3buHsiz0Akn0mZkzex+
lo5QOHZEQOUIpJys/6ira7fAbYDXDgUtUrj4tzRnqg4Q8H6WyIe+Vfb4CgQQ3PVdmXwUIflvD29r
w01BSqrqa1wDIL/KjbEoWQ+N6esHIFCTrPYdmaOVFYGhjE2TGyUNXo/iIqi50DqOnW+72NNu5+Ht
yJVHc9rmgdEOKEDQkDSygYQiNbGNQXxewAfd/ox9RzFxtHzYTSi+ECgx8aRylgRNg+HvJInmXbhQ
mqd56WS4wZeqg8mk1Srd77Iq0ow9MWQSxulr6vfyLIyZBaybnbGV4L4uCIrt2KyWgWux/gyLglKK
Q36jROFC/iq7j+fDbHT7YqlYnq7U0gcIkiyf0MsPVk8YVSuLbzYbvrjbCvaEaZATQQVy/ofdfsGD
bWZA2902B5hnqTFMiTt0zHkKiwyATwdSDKtkyc/JvQnHidMsQaydmCmEvitsRsDVT+HIKgA/SZVu
Pi6S93io97aREXNbtzjMc7eaWRL2LzMyJo+SMp6I8lXphxGp311dnCNRXsLuvGJ8PYUpptdiAHcA
zmVLAzoWii8xNwjrfnj50iznzMlXk2yvMr0wQ9f4LhZbsrRq8cRyoGHBGBv1FIp9uEiD1HQg+zuE
1euhSdHwLioAk/tXmm02Qy/tZqjaEi5jIbR7jj+80Zintiv7LnkR9/q85S/ENPiO+gyeo3vnI8Ta
DkiHkNo1HqSPitdatu/739/mAmyaaORuLmMP8zIj3QxdQDKG5Uk5EHzYunrGN/Ka0w3JxrVUvHBO
rW2bjvZ4/c2eO4znKBz12ndqX3G4LI0/sKOaX5HFigA7l+CpPZpldut8gyQakoaxjwe1hcCqocYb
nAacBtmOlH/5rkpvM5CykUXt0OZ9jF8zw8Gzi6b/EEVasiRui7LLvC/0UJ6uMHUSdGvNTnKfntsR
JFAZk4QsnmF+kdxneDltPRYpnMfI2UT667a2XRt6KkucbrRlP6+dgtr+y74AmqJW7p2dMUBWTJR5
U8V7vo0GMVGe5lPTD29gx8snM/2Ecf+Xqy0tdiVDaJve3lWs23nbrN1957ALvgvFHjoUrlQLjC5V
2kUBWJ/gHVA8FNuwQnoAY3H3p7ZLwA6MtYB745Rxc6EnLBt9QG56sl5UQongF7dqAbyAQc8ioVwI
Lczsx3hC7eA/+3koFDoYdGZUOiQt0kwmQc/4QekaEJC+AqFO/PFNyGZ1fq36x5Hd+x3q2dJGN8Di
NSy7ksRGmSgpV/osirUM/PMEr97w7WAaJp6GEFzKyMPKpAi6fr7QqKZ83RNyYytz1qcBQRK7ZfqC
xmffJ6dlnR8Thh4QnT+b8EFKj2CjaPi3/UfTBx1k9mlSfSFAW1ZGC2xgqvQJrZRlWAAPifeTY3IL
B16mcioGZLTcOSK4DWOpQTvio2K8/dZJ9PHndIsixojmHyB1sSexbJ/hRAyq2RpFl9SK9usIlU7H
hDIkuKKNn5Zesn6EKLmy2KIUlOD2EsLyEq4zH4B6w3RBwOMnbNDtMKwUhbTPjMQhjzFRdHo1Mz/+
9WonrfZfDPrAVSqzvJ0/e9/x29aSH0yVJV9FNI38js+sso7njxGBRsNdVc7CpHTZnl63hHvmj1a+
r4C/uV66/4LIQsjFNTzrFIr6XhU+jKtD17vGX7Aqb5Dsgx33CS/CgCejcuWcM//MYU0lj5ADKZpC
XkklJZtEZXV0DYN7uTBqNaAet7Bg9+WaydMmIcccEQrRIqPct9nGVLJai20OYudKphKMIx6dDqxk
TlqhCROVl4tPp9IfWaxApaLopU6R660AnWy4dLVwdcZxVUdVslPO88zcHLMvC7qHEFf8tBldaN+O
ZIkagC3UMmy4CEO3mQY8kE8A5Tu1cSRgIuETTPKfo3ZdoN4Q6wDAo5t7xOwFBfCoxP96Kds2auC4
sdzhiHwnPnTaznvytEr2jECXztfIegfzIR2FkD3qtXnAWK90n3WYBLGtsfq58er9Jiyn4o+OR4KV
vvAPHs7OifH3hCy2vVWhRyZc40hsL6a7PYnzMmS3NJyc8tqYE7F2TgRXiAhkYX3Bar0+2LlSvwsv
og2eH4hALoGQfc+4F192i9UQDyEiEXlE60DRIBeEVYUBj5VP+blfRtPQO5WGwZ1ePVO/S/njLJUS
3us1/AaXyBEOlfcMAQwHmLjp3WZ72F1nCPAXxNpNw3AYS4g/MVt4VYxmw175lvb6tKAzxikQael3
2IcneKVy0tCLvFbFcoqAIDI8bN3dcbyT0nKd3ynrjk3iiu1pZsBn7Ns20MK1TT6wvmoj/r6bgiAY
iNQhsMh93Zwy1gegB/EqjgD5X5li13LBFIwEmgqOShCm5glsVQaaqU6R1utVNeRqsK+Fp8SYjKKQ
OOjNUqpH4lfhFnrAymafJnTcv1Slve6S7+lObc6/n/i3xygMdyzcOkvTivrmROsDd+qDlfIetPQk
CmH2x2Q6s3w/rdmYC/6gASm/i3iYMrf5GXWkK4+tb2D6Hf1YjCc8tYZMfGjDTQNcG/jbYTiMdNaK
2fCMzEPkabf0PFDuTPqeohhv//zK8NmDOJkxfcRK9XRpF0E/pngWWzOfvjYba6kAxAcvFuamrriC
grcXiDH+B9QbNiXr7RbOEj4qUlZUOu638rHqDl6GdY/hlhgWoEwY89p+4pyS49v3yoUfeU0uhWi5
LPqOaS2TSnc0MSMA+Rg4ez8Zj8Y7QR4QqI0sin5HvrITBVl2PiNf5HeqqNVUDnfTI+W5wN7gpAV5
C1h0R5oQyaLGirL9iiv09Mxak/8QYP5QmENBWv3cgOYVii6mpwth8reg3/M7UP4prlt6UIek1MVU
3o3I0kTKXv19vA34Ctez+o1r0DzzciRla2CKzD2hl1MFXf9Z/j2wiEw8zPbgvz5GOOipB+mN8Te/
tugZYFddmCVTcPQzGx+Ch0c9H3DeFh26kQC7Vb5BUxfn91rgTwZZbrnEmaRY5dIIcYTM1tOa3/RK
brQBXJ0CnMk9VkjE5zWWxAqGR20r7+rY4VnBvPiN6R13Vr6Sg6pon0HXd/sSKNQ9QKiOhLSFeVK+
AzIm40yMu3A9YvCQlONi46U+hT7kspMuGw9U6gd/HBfybgES0GEl+QUmOJZdwkANqprPfBhVsy+h
MWjKiZAExxAQtg/v4RsVgpa+eQWVHz/c2+tRG/IptFSJJEbgvUDybco54m7ahckvnDO4QNA0P4qM
0dyCK2ED4NoFbHJqPPq+Ojbqjdk9MltuC7AlHblVuvORUoQgQM6CDzJcDdRBWCF1DPIbwd3wOxX4
X/3zPtewsSxzu8wBQUzaxG4qKfvFBt3D/NnWANJn4NlAy8bhadbHAE6xaDIyTX70xEWAG0adzHXh
yYdpcV6Nfc2oWLhC1GkCMtLVWGxSRNMUp/WaGkPctKYdKrIHudqNEWHEHXYyA0WthrBBXWSR5KKw
AT4lIEuYZJNJoGIlDm2lpjemIHAZt9VhNG7fobQjdtz1XEeZ+jA+sgg/lIy9e0DUVsz6WHBx4ZlI
EghZl3SG9DcOu1tchwvhT3LhBvG4hZPnboxkMi63f7cJz8lzSNyuflvf7jZImFJK4jOr6gEa8OL3
xomHjONKemDq8524N49+h5R+xR1ilEgh6uXQbRx3HdIPZwUpmo1UW6w7LpX4IKHKMXYKS3aJ5/k1
Ydjd5q/zeuX3DkdaL1t62ztB1Fd3rB+mFavmSPVHiZ2oEvzPtT8wvk0gDhVRn2uYcNGf8crtCRdB
BgI3WROpHDLFnReSHV4MWtadH73ES7HrUB9USWWWYPLnVOQPHfeTyP6VdLtSJJplBOxdLJbbZvMb
QDeg+MzD0T4kT8mY5R9c/l4+W/oqiMeJC/0xVNbKLerZiNy8pz65XBO5z4LXZBQKVhref+9YgJCU
GeTqRidHb3AKVCQbMNwtHTYOL2fdLxKry0HXHqOguIz5MjAEWl7/jj6d/B/2lt+8XiiLG4XxMgK6
hbwuiESqM0yt7HcHxDWM+UyEV9woHGEBjHWYRJcB1PNaDvMN9wkf5O0xcRPAqQXpfu/NoKIUTWhz
MewHqmf/7BIX5b9mhzdbnvaAijiXXglyuZowQrYTweHTYVbFeSPy9vgKeT/0QOop7GKefeYa+Unx
f08fSZGjBCnPkJkz4D9KsHIxkD1iNbXhgFucsD9RUZ1/spzj1NEYNCUeWuFr+xYmHXNhFQMtaDZI
uhZHP9dUQGf7W6Rpm7NleFx6hWkQUICqkW+zer6OmPZQ5FncI7uC1b7QwQSpuZybR7gNPp882TBH
J/LWMJnOVEzJBJ3gAujFBPPx2imYozeE8tEXLTxohV+n0OMgZ9GbQGoQbMeYugY8CxF8aRH9jC7J
PFeuFzIPAl9MSAnuqu8hTMJikeV9Yqlqc7AvIxpXY3H8v81IgbBFZ1poKdzfjWAV+KMqVuDKGCYZ
GETie6DMHkKFvUdd06+lw99BBwlqiQ6BOEziWwwy+mP5fnFMasdmUMxtwQfUe3COMYb0f7yme4fw
b7hoqNUY4OQvIF49uttyB5oBuxbQe6LZ9tmEVuPmHTDqLBH4fnoR0KvK8d77P0RrEu+hmFiEcSV1
83Al/5OJQE8Loqbvqb1i6AopWNSNFcCfXF8GQWxZFcjIuebnYuNFubS4VlqTNyvxGTpYUnWcR2C7
wTCuu8lA0YGXcXIU4QVoCJ4vgt0H5hV0KGUgHCv4j9SbFkH5qZZQVQdy9HpJ4piotKjvIPPPmpNc
p7bD71BWkR/Wtc7YWZWqSokp4QlaII8JwOfZOSnis2+LT+JaTyjQk3mLFf5l/xyMeduVJ66PM09p
YYP/xctD8DACz5SfR0xZiE/BMRafRhh7z9EMrC+lE8mtUpGv50d1rLYNEWu/dmV9rt88EFuwUdAH
NrJIZmuoiW9Ok89tnUQ4FUmuw/Xpr1X+Uy2EWUgUyOljeY/5Y91WYGTYxrxM4sLdRm4U1RPYgysd
hiN8ZUC8GmsUmFtWhSpbXNzGxCoUi+RVaWaDyKFrriee5ILZGu81s56KjVR0N4fZMr/h/Jh57aJQ
XV8QTMLFrZAiqaDmIDovsNnyOUCFnrwU4A+s7uqodJT0zNlxeLruqummBC3veGbC+eX8X2XloH/3
lCUtO7jgCyUMRrERG9unAaEPC22Q3jkFhgvVH3nDfsRrKaiUi2rPf3S2LSnXwO8S3XrJ7CEvWXJs
RMrCN+dWn4rIAMdzH3t+1Y5QfdUIefleEkblFrgYtgEK2naHaQwhj+gE4iA65wqLXOHMVf9gAMiP
C9CJqWxsxLJT6PuOMpkl/mNgb14RWZumKyMbv7ub/9BR7dV8I895rr9ECvgS8vkjhtRgPe3UTwQS
+hgEdyYXtgISNYBbfdiAMv3lofAjGEhXu3jclFan4+bDWFhmy1wp6ypM23Vef2GJqBxI1kWfFJCt
ff9JDdvjF3R+y2sATmp8kWYhHUfmc2v1+yvv1un/dXD9WjMBfQuAZqK/aiGfobgvNH6ZiHin5gUC
BlL23ABTlahlb1cUG3CafDixB/Bcs0RiWvpwFdYird6TYmDk43MuPjxQwGQz36Ko88LplfqZpLmJ
0uHp1TY3n2V99SoLpl4qBTurLmwMQN9rOpEUlo8F3GBvKxh2OtimVqjEbSceRIriKl+HM174xKIY
BuhL0Z2iO2riwMYMTWPYz0bcU1RlspTFrCU59R0VGa4Yo5SdYxO7an16vxLSqlgOcfGANuVIDF0j
eqb50m72RyIiS2Dn9qfuQE6bJHJvSVD6P0TD5DDlwASyRtYvNh9x17mjtkR30N69P4v+dq4PfILs
UKkALz+SWcQZYBEr2HLpi5ZYNH4VNCY1ZzuTESP7ZDEnFmfw4iv7z+xuAa+jVxOMWZ0r+lPGykwR
fKk8HbX928qswN5HA19DB/DWLPrXSyYF1AEteDAi9gaQOXiE3zXCOCWlAEX+fbTj1cDwUYwy4ywi
vfse1zD8nQsOL0/4N9IX4KxCkAOsmdRvsp0mOVwo9hLE1kxCk1Df2aY4kRgauhEksJCKmXA38M4H
lpEi4n17tPYGP26XZLVctEYFD9a/GwRnn+K1WehaiBUesjgjP7DqHpwYNwitddBzs6mhyDOL6m1E
2Yvy3iuy8vpbun9rIpRV0VyRIdFxONV54rCLzDz8Riunjk6UA2xBge6cb3NUkyMb+z2efUdjhIZI
2AUaJWJpq/wIzFdWhEc79RIWOOI1TmUOYjGvjSLMX/D7p+8H2eMIJuP+lukACP7Ssfzz+x9md0t5
hSztsqqFxJTs0qNgj6ALYeD65mw9UdTpBnmUHhKxcxWvnq3TsHOVhcQCDgXaGOmkKMDQMm4/riCQ
wGu7xTbyCLZQTfafM/8BQTa9noC9/O3UUxmcgftrLqePHsY17m7aujeWxB/BT6fz1us1hzDjm8b9
MqAcRq3y6J1h1+lEnwAJkivlSma+P98AGtijsbulYijLDMC1uKzQCokI3OsGKWNW5BvIpcR58Wp4
KAo8hkkFirAuf//SslnA+iFacpoZwkaGRRXkjwFwEZ0INOjlyOT5uhS0XufBceSZwIL40JW+boEF
eCiaD+1iur9PWOHkMK7Z3mgcqaith5Cyweh22M8KhylW1uHQFOdEpLqmCM7PPRbK/8kRlFf5JriS
1nrCt5nsnf7xa1e05MCbhCPK37dXXjZx9AAU7Qb79cYQ+Lk+TjAbmF0U01R3FnGkWMTtUHg7vh3c
leyfPseCyQr5hr7jxfsJVPlw5aQrtpKrxyO5/Gof6TgFX67qy02liKPKghUR/53xHKTEY/gYEKR3
KSSqA65wSP8A8HFyiwv2s0qUFddIQyHZ970iV9a6QaJBtbArSodECA5x/3dHu/4NqLbcd5uS4SaP
OMNsyxN4VC26f47gikc/UkdYg23b43WfJ+oefPXu5Z2buOH0wqW8cKLQgDGfzgBXRr6YB23Nb3ZN
ODzaZ5W0jpnVJo3FS7RAoVnpxaCNl/KjvDMpGMUCnZ1pKenawIydmduqViU/ODgp9Z8b2E0tAT3i
wQbOGOENfS2dUGY3mEvxlUa39typUVdiongTf4a/00XhmrOBQklZ8s94gKc5dcpuOZXAm8RvgbqM
Dx0Mm0BUJaUlEfyQTSg6BzPohl7GtriD9Rww63IaFIz4EnoR6IU8MWp05PVmkQNemzHLrOJAzQ8v
kllS2+XZ1Ny73sOpPlBqIsu+gfRSPJBsSiIVQye7pHIgJBrSJfQum0NJRBwZbYS6yA3fLjWWvshS
3iCNftGFtDP2VKT/XPTXVnCJk9rHRGNd425sXODP5eZAIUvHD4A9QQQT6VOx3GfwoK+Y0HBRXScl
DRvBBanS3fZPO9elIoPSH0+B7uIVDw5RdVeMi6kvOqcCJLS/RdlPsLGPjoQDTJXdNYCJa+lyL9TC
bgDLNbXcfbkDEc3SbZ5bynuAtSfNfv9zHwBGANvLX78gSRqpLL61hYlEMOkvlacM0k6jfuuXkf5H
EaLD4VIGfj6ocduDwmwQqpHdaSYQE5G78Dhn0LjTqGRW0joNg4O8aQ9W+eLPZyntJxE3hGsZDtXW
zc7UFDQn5sjeMaiNSXKDOoyktsIqgK3cBNrOa9m7O4X4p60283rzr5pkLv7EMVi2sXYhr5fgddSG
H0ystiPh+Y+zLPhry+gY/nTl+/c4I0BsIhEhtnInxf9aNArFCjYt4Jokezi06kzGs145dYO5zIgv
PKFyM6Y3Fq12VqzN9qjWh+k29hseiphtYtfIRVxYMMA5MQTHaXVJCe2p7wSeq5O2jA7FJ+rUMRbc
XcvQMStA06eFAI2MYIPuc1KpT5TqbzJRLSqWzJaLAFGfc0X/86NsT1XM39d0bhi25LOY4zVOTlZY
g+LgITqOFJp4IegWTEC3NHg20luCGD+VcRTD0mDFVRT2vpH+6b5TjjhtvwEc+FVrmqTIxvzjqsdv
YrbALMfP4K1iChcM1Fqb2mVb5gAyeEe+8/RHP0kM5/E81QD7VmMTabTRMMW/Nt3a3/ePQMlWl93S
tWumiuyYTjAjGSGSjEizzGKLDSYPLwOmPxd+fgaTsS1D4KxG55rBpZE6UCrO2eCI8DVA5oki2FR+
l5cZQehHfAE6ChyxBxqQEHS724PqtJT3DblJGI2Y/06y1EzAkc/A06SIRFeSV3rwq7vkpIITG7cA
N5HYWEOgsc1XMWFoQ7GBzwS4VyqdamiMQIS8qjS5DkxELBjonhxhWw1SOCY1Pv9mkbN1A30CG6iC
CC976W15yo1ZlmyqDEWmA51mf7GJSJ9AMLdIGLdMU7hEdMPUlZGj502l7g0V4Yo8DDQl92XN0TTB
hn4IoAb1nVj8XaNyCpdnV+XxaUOOD+hj8yqm1PeeRnEwYjFqrDyThLgEmiiNTbXPZL6D2Pk34b2g
cll8v1adB6+wC948tyQopHlSvM9VxGexRzmnxeH5W8hBvaNBBZz0AqL2aVrg/N13mximUdmki7o2
xYt+WH5Vht8S8B6WhOCQ5mmzDqJz8cOL1q7P2ca6wzKcNvyMTezUg8dYy6KQcf851bxgDXvucJDz
BiBFiw8YkjVS09moc5ibWtjKjAGoF/uDRk497G4QfQ3XSgSzxVm2ux3/LjYqR7BC/XUhcRJz8e5N
uRfBKVXeEwivNPeo9dd00Hjl0iwLb1xy/ni6Fk7czU2NJIAwV66avqWMzi4Kbcua5YcCzVVrJ9+n
83U7NUjognvxPKMH2mwquLuxW4JbGy+2M8ZDGfE70shNCH6dhyICi/S6JHzMT+yZhJy0cjm4qrqv
n5qmZHJst2nnmo+pkBKysohRh41m8vAx/T4jmSXUpu6eQQMCQfHfshQHYQaUIgyn5wazgMYov5PO
hgHGjnGAGvMLBYKlXfqODxH2W3A/cy86VHomPgreK0hsM0snsFwRikRBIkCca7mGwzYps03syDgd
61dgcFtH8Qr6NApLy6TiyBx0M4lwA8gOcWlK12YKiTOzn332Eyts3wyP6AxDdTQTSmrsImclMvty
91lix3+3bs6yg14TtVQ6fHWFawpsSlM/L1Bcf1JLZSr8EIKH9/HUmok/UPjJD2LE0zTnGyZ6OR7k
UF0cYVSSmxnnxeMjQ74WHdce7RN68+38PC0D4QTkIKP3qmOIKVXY0eaDcIRE/9MM3OTT0oBnXAuu
JCnavYzMYA86RjKGjdIFrm0pM+BOkNxb5Zexa527vxqQcJ/L7VzUoorvOKIY8rJJoixAPcOCLFkV
fZhBHkfxbfT+YE+EQTSKu9rVAH2VOLdYtvKbmY2lXBAbB87M0qPbQu3esoqClc8LYth7PH9+E2NS
BIvdkTYRq28og5rFV2Mi4xAZhIEXg3ct6odkUOCLI61RMrLgYEWkIklDHw/1KbwXF7gYhmHkajZq
mB6TFClIqT23qHH13V2WlnxL4/zS13CRAaWOYuRLwhXaNnrkq6ty6DwfQs4xzYUW8h9uyg57ZIMW
moX0QcQc+AGdoU2gbP14pI4Yzao5UMkdywi412dR3pG1bvvd5ejX8rAPFPJKvgQKQmDWuDpQZ/rK
d7YOtxJW1+LgyA1zBIraAahU4JjyBOJABhiIf1bFZ3Z/j3xtaqsxykB4VlllbB9dICk7b/vuh5up
vKfpky5+7h6VRoKC6WBOFP7W2Qvxh6OetJaSAzMsq9Shxx+2YIirR/4rx9ZCydAEG8Bi462FblXa
2lVcz15TvNowSKQwEK/8WxLdRO6CHH8nEOtHanzsxrbfdYf4AUZOvhp9oxdGzZmcOQNeH2NaXsWd
sQHO8x9RyjiIBCGqNPKWTb4ooJioplxQOqn0HdYppkdQN8Gd/gI1uEiS1jrS7xwqV8uzuZsc5JuH
N2KQ/dT4iRZZ02uurdDZIVT/PDY3yQHbaAtm4vS/mXWuZV8b/iJQVhSyoz1f3NglID8pfStW6LET
9KQxqIL88ikEV2KTTlxCdTK05Z2kSO69pU2UYX7h+q+iWEh3kggXyEuESjAojo8T52lkOV3tSN92
dVmSmKfCkknwW7+i2Dk9gf/eHMKu/U0RqOB4KHZ36ShaFfABZ9O9lCiDEZYiUEL5M5M8mBaRviab
BlbqfArpqf7g2E6BQqiQwAp3jAVT56ZAi1NKyg9DWv51uBpjpw6dLCHtaZkBQ453w1B6FCzMJhOA
T+rHYSJ1khcjII/jCarj0gWiFXbLwlD2YNweSeX8E56FO/EB1FC0yVGSob0T2Byupmh+zq+wWHDU
xaaSqTZLSVWNy0ASr8+oolnlSzKVF3wNATDeEhaZbZ5qLxauZyt1DjHg69Otvv1NpsBz7nlh4eHo
/+iOD0si8K147zH4RgfhwVK/5GeEWB34TFy9hdhBzjXTJQT4vHIQiSWsgBbJ022BCuBgf1pXAbhu
vXJVA3vCorRu5+H1m43VtiCUW6oyjPNfPFhiMIP9o0MuJaGsKBXdWCATq1Yl2FcY6ORFuEmWr1xW
eh623djEY3++/t2fk7qIqTpgfC/tDaOMjcSC2TgkoCu5gDV8ATY9dOuTlFBQsSeH7dpPdx60EoOy
z4IQIX1vsOX4bnojX8YTdJC+TdL4HpDeGPNO9+SJLFTZPBPyVcXpu2CKZfE32cyRDXAm/CL1toVE
CWhOdJATGKrAR6AX5GY2DOYYGpqG0pBPofZtTIW8owU4CIzvEzbG2F9GZauHRSAW7TAEcN4eGInY
sHWbcnzzeZ/nwSMm1e/5FKyoOTBswFWOf+WqnQwuNlmW9dna/KFMZyJT5Mv9F1jQSOoYwLND+H+B
7lvxqw8ZegeBJ+hdyWb2zqtogfn/PJJcgoo+6thkATOL+PSp88WYpOCevFhXHkJkJIEMACKfnCXL
uGlYNDf0FTHwg5HyibYqd9L4zIjhvAPJl9t7I1glOU8/+ZmGn0j9en6Zp2sbkcusuwykCwxgiCPS
1o2dJJ7DFUwh35HTIHcq6X7lMzRksr9LbjhIi9nell7doupKq9r8Sx1PWV8gdxjqNLU0hyFeBw16
/902DvBPic0Mez/qyx6sV5XHbxBl83Db8BY5bLB505nkCs4Ogm60JaqHgEIJFnhSulqPY4Y6kvPx
F+9QtRUkoKPng7OMXH7cC22Oh12vrEam/VoRDT3qstJJA9EX0nwkYQCVpJt7NMUVEKKktZ9qb445
TummkK7Yndw7K3UlP5BRZ9nqfRZyiaAX28Sd+OPQnala5iv4/XNhzmDyvgMqz98LTIyd3eTHGln7
3NFv2pJ80zep/lDnFkyZchJppPR4P2+0AWbstnlIzd28WnbGfXb8o5noP5jN5FeSyyyjAruyMAY+
9uX2SqXKFukzQqRDgbPh/Glahy5mRcAOOPh1yZyatOINDtgrtKLNEpncVjjs045dSffSS2dx7Wye
K1vYOvhMouqNQ4DGd9UlZNUI83wqPyOTubEzL53euTGO84oD1lFr/owQ8A8EMX8tyvct8EN4LvgS
/NEv938HRlizR3YZQeRXTEGihZfgVhlnczbKUnSVqfaetrqOuSINVrX3NoLsMqxP86oMJbNfidNL
EVs8UImU3Y+T4j7gFnIdr+4D9inhOlW6htM17Zgko5tHNcTR69E3MdptLDDsJrQawuesfhz6bWAI
rJ5r0o4iJRw3ASPNZI7gGX9rw4ruLpMiLU9dGNTMsmuBB9jdvcBPNpq0rEQ07fFuJo4eVci5cFfL
ecAxKua2g2Nvq5sBHJthaD1L3ri31teUamAzAXfZR9Hz3dh+JQN/vkfj19CnnSFUPEzitZa4JUJC
hkAaye7xkE05sP/OI6sAnq8f5ccw/AqnPp2xDBb4hZIbJtuL3UQMxemnsTQJnYGkYvsR2u/YlM4N
QmnuUYSm4h2rzfaWUeO81j2B1GzEyJ0kXbBlBciuhnlewI4ZtxKuc8Kje+bpAhigAlyxCqz9AcS2
8aArIGpLMkeyFbJEQCGRRTK06vmJc8Sb0as1NNvXk5dKAgOOimRav5wW0WOWs1VrRSzyRmrr2esX
ssuQYdeJoBW7+PH2QdQ7vfwCK0xS5/Q0eUMM/9J0tUlJp+wgzlcP4KxZ80irgGpiYHBGtVE4hylG
6t2ppLuOasdDypsWWb8D8sfr7F6ywMjcp1qOTLxqv1DVfJPLlyzPw3qA6cfziUGmfpfWVcRmHAhz
PX6hjCOoXc+pzDcw6QflM4lzV25ehN7b/6dB7/n1+25peZeGZ2VfOxAp/VYOICIW4RuQX9OPkp/2
WpUC2D9UVkmQhbQlka8B/X+Wz1sV1HitoYDcx4ZDb61uXEJTYtlDDK7xWuplzfhQu4pjZiCdxPWl
OkF4H3U610ehupGHzSXNTXUQpsriobutBly3Pje2b9vQB0tXkdSusR2zzxJ+kdoOhRK8qHFIzGA5
rSCKhgbtLpHhNrz6y+5Zk4Nvkj8gNDWXuTg3DU2CTAeuTvdE3IA/FgF3dQkhow1yg7sGu91zMd+Y
UE/bDU3rt23AxMutzW9qKQ/02s/+J1bRhJuyeuZ/KwlkFtgYwuRLZRDd0p5cv7s+y1H1cT+Qgf22
KErz90aQB4Qmba7sLLjHXi7zYGlscZRzi1oBui00VZ9dZ5oLDmc5/H+CfAcFxR+j0ba161+6Ce2r
P2z+e9StuEcRLsE+WPL8uxbgd9HG/LusaWWDtdc6mHWtxjJzfFLLp0J50tOC40B3zSRXWk8QDiS0
R5+GxGcYgbKulh0+b/+PNpDhEfwB0oVSdN8gdSPNBCbAXqWzcyElKeCSV8oyaR4nfIovVdaOmM6z
UaDysh6B3kRgasxwtJ0AUxuCt5RYGKjG6d3YydB/tu7oeTIScXiEb1U0VoJ9xly/Yh+BmbScHQbS
rj7ztQsJeTcSTfXVA0jgKQF7gG0EHbWI+nhh2lhCemaruRScuDs8AR8vgvDcraw6GkdeNpKkc0+c
N09fbXdJEM6us3wmpXuVMJO62ioFNrbrSmXkWcp3CJOPWfx7/HxJDJuy68gT94dRZOwzH5zRnagR
GIj/b4ZXJdUaQq/QTpont998jjOrS5nQLSN6kXQeaiQpNvwDNX+SAvdbLPnE9SVB5D/OkoFuDZq6
y9/NKZ1p2BHgTNRStb3ORxiSPXAmJ3MH671iWI5ty7JhYOJkCkSWDvgH2/rSUaiC05IiZ7gKUfH2
7it0XjRmP/cRKXhRP/OJsrnGlKJ9wNcCJkF5LeDRCRe5GeB6jBhq3nIbjNv0rl6boHvH3Op5w2vi
cGYEjtX83vCYg5U3pXqIEa3hv3veGosmjH+NBoSsYwuTUrzFmZRzDN+zpagQNHTZhMD+avvWRFNp
sHLBjzABw7IK3XouXcwXk4Yj5/h5FWPfhnuuhX2LGoPWtXbQ108PqLrkxopg2xvR/0ptQLHwv2qW
jqG3rqTw+W8zhfZUrE6LItPWmceqNDxqiF03gUm+ZpZfoxRsADJ6P5Im2yp/u1UQJYKG3rLD+tEX
GUAS1oM3P+qzPTfdx2sL2l0BLuwYEMDEwz3dNVcWEKMJ4BjB1hyij6Wev/MnF4OMGGtfcsGWICcT
/nEiAJzxWtLa3DBaiK0w2SJjrvtpea63QfigiSXgVeCnuES4/HnY/zN3ShEsL2foCauL2TIQb65Q
5EkWxzLH6OyGYImsr9Yfk5gVnwHbNMDc2oQPoFVgghPcmHE/ufSrPS460FibYF4R5o97tSrdLw/M
JMj/69xqdxAdKsoLXhmmZaLCQkANPtL06TzfMW0RoONikkAL8VQDwhkJkvtNz5tewUCU2NurCcnS
iTBbj4fBRfuoDCdJtBY+8Y/tyWyYc6dIWI/Hac+6YokMP2coHMqawG7pDU7y+8HTUIOa6aoK+qh6
YQUbJ6cPLNuFHj1bION923keX/uKi6EvUi2kS+YTDBu7tNa2mTVEWyHwW4TnBB4OEQiULaZMoe1A
uPs20pS2ER9MkEiSINAAQlnWzMlxxLt2o8LFuOWQyobuCkGQLGZvsdRl/OsDdPeaedwk6YyPUJlZ
3vQ7Lb0E9iEtXWvPbzTUOL3e3MVdOLdjdBOYPPtmZU3hv8DRyZuYzVR6AL5nRC83WNZUz7iRVsAI
W7icQHDfa7doz+7Sjz4iHjfnVK0UKFFtewJAKYR034PiShHdNT7Uq19SV2hNuKYW7o0hDeG/X9DG
EVytqpWsXlM4MY7SC9LclY+0QbQzD/ibHSWzblfGHSxJTipZSLJgFHO2GPNW/SGJom848XiQuIU4
hb3xp3r/XihNnQ7O4ylZjVJrcC5T00UWbc8DDbVNpPATBbv+ke8sejvgijw6nA7AjY2Krv3mKntF
qkxCqb5mg+rnGl9XJQUTRXMukusEpEfO4+u17YXy4JtgNBpKPfDEtfwx1jJfKX0b2nCivobAohwJ
COIS78PabDA3WsUWAfLJ5S469/ZqUCdjCooz2IIPjX5W3V8dUCbY9603zqKINpmbfGLqcQ71nPAs
YQHOTZ59cW0GQRpAntz42tyEDxqPQbbbEO/WhViWdPaEpvvLJO9hMtaZiOZoFS814/QKwCwXXPq3
6eS/cINMqW4fBvEi2IwhCWpjih9akIUX3HatJ5YAFj7Kz+swV2KENvRwll5ImJGmVtke59X3L8NJ
jCQNY2GchGUVANqQ0vkgCe9nCsF9dC3aOMsrdkpuMaQjqWH1TJ7pSMXVCoewy2XvIcZ0hg1UCTpX
L3ExNqHWJCHVDy/QL0FmGrICcf/1K94W791mix/W3L2BHsYCM0LXFRmudaLC4DkUfwpKUYNCmZYF
ehr4faK9ghCikNpx5cK3pKRxr7rEOpXknXJGhCNudDKPV+O8PAwXy8u0wALJtIDvRWd0XEaxUSlW
1qTgj5jRQXbn9BMPVjJTLIuMTtBzFIBuYY6SsleuG1nEeRgYaOSGP4iWBzhOFVdBatRIsGyq5acm
rEXI85EU4Oma/nNxdbiWYRQsKMdmmf4NNM2L85TX+TZGf3QUo2ABBsbZ2B5T1ShQz95FbcEAVqD9
vRhCZwlqDbrsrm6ScvNy0CDa4eutpVgWbQo4Z3hXWWZ8yOzB+fiNOLEPpCuodbJPkXnspOQ7U1wH
lQYTU1MnK4Ur55c9/1IYgqCwN4rG5lg68IKl20VPNSYeKwBgQniyRo7miRVlYSLBfQvKXxNJXXGD
OcaVafiP9qnLsQRqBHuiw0zYrCh2pWFCFoTqs6Ofjclgp1edyT7zljM3bDTZNOkIO/Fga5/DXSTm
tbCRC65GMeN94xIqhp/nIkRvGHYXx9ym0xsyEYfvmf2CMwnvI0HRndQSKjlL+RZOj+eJN9bQXPQj
c1vJxcMSHEqesp+TSKQK9SpYDge5v4NagJAzInTvSgiQghr4nfd0kb5JeziKHONN93kvHXnruOzZ
eVcqo1mHOAmMStUzRpT5/9+ozYbQ1u0Zm1BWosXN/vIAGRX/NaJIWhGDWIm1/5aESD8WfFZ6IaZn
W2MnY10Cmnbt1/KMhvMjmlJVSefqm35L61hdSMHbli+u7bTFUxB+qD+u8IL3B0gP6sa47QVAuktF
HoxmdNSv6CSoFZck3zrpJT+MNU5aiWzVrVfUqLcsK2qtdm4VLsjZYWe/rpx7TADOk6GyevkZqeZl
hcZcFDhJBlEYs9tXI6dA3nEuccH8mYTM1Uo3ZBXmayiAUh2XH2Lw3/g7YNmlO4Uhf/9O8tMVoDpw
rHIfBz9vPKkaj4OsqyT+buZfbt6mh0snwW4yrSny2t5pRDn8yYuwnrXWfkKTIErAx8ZucbfEJPyL
b75h0NvaPtRj2iU3RsSVabdp6STi0TwntqqWmVc23CIKxHTIUkc1wD8qsjFEa1TyE9ljN1uTTCL4
7valBvAn7g38x8jsJgRfRJcWLOHkqU8D+76o0sqtRCvKMTU7YIQm5yLbbuPh1LL+WJT+5YK+eg3r
/slBEsB8Xpv/64rt5qVk5tNEc44MgFFkAkpOymJO63UilxkAoWDoCLcA5h1XTsN6CxJQEG4I7UQq
AUxoMkIWmsrLvFC/DRrV8TPyvz/9VoS/WIdDYLMvs4nX/Guw8XxKma6231T6Wl8DdQqgclPFcZIS
DTrAZhvWFdHcPUjDzhZTDPX4Zg9vkpOGHwxPHL07YfPauuBVK+ncg6uHp4HZvxfAa29t0LzAcddj
MNAQd0dtm/RMaQwLQBYrjC1VFTA5rqIuM8SW0ENu6/MeVXFo5qC1zzq+opyY/hffVAl3U5fFdHXs
lj9nEYpVNlBCslZA/hEhxCqEqRwb8OPeWLjsA7Vsi0E6mWOeu35UX2bxVQ4U7Cyd9z5XMCUH8UYf
XPFPALIboI4ZAFra7lY+gmDk956jPvP3E8+HY0v1fBpEIDVk65JX5/isQscyR1UFy0+zYpkHRFCP
bSCeyw56/ij3jbClbOwW8S/+fnOj6/IKAada9aORO9eB/M+a03HLrgFR+mIU6GUXttcYkr2dQMGR
WWGVILfSRaAYZojIyktUFXSuSQJjMLIyvKTSvXryyGtEbSX07vDnHmTihS4R6hjHCRJCR427Huc8
J1kPVgxY76G2hdhd8kLCTjJtu0gBAVJfrkygdN3QeSPjS8Mdzm2Jq+Wyr5jI1r5mQ7bCVTYF6Fi1
f/6DB8k7Xn1qKNhdFaQvS8MbgSa1czh62wgqd36ZtvjT8F+HTmPpcFSpk3DJG4xI2q38LVfp9rvG
xMG2FSz3B9j5LWZ//FSC6ubFLnQYOpIKP99Krs/sGnuxWXY6jiOTy0VeM26ODy/2KefV0v8jsRSE
4Ppx8RE0EkSlY7L7C6EAxn4qmu6+snRveB1vDgNjbgdbVLhE7qbI57GN/i0jniQ5d4loqjWYIn7R
62vfuQNz5+bRDODEFNNXVeJ5NE9Mtb7ncfNLZY7cNRik9bavatg2Prs2yRX0flzGw/aq1zwZLPmR
Pwm25ZAEstN/jv7hEiNdElBFn/H27gyj4lC7hhunX0NBLtIkbENeLeYJyW4c93nDH3/zaD3KkkuZ
/ZrMIgcYESBV9A1/bmrj/zwfk4S+dZx0Rk2sWIKvRZnkHwWNbpn/vF5aua4wcH10mQODVGh4SU3F
G9d6/I1m3Pa1CeEoEgvIeK/JGv8B+t8wy3wO925h4chYEVM+TpIC6lmuLtjtIK6H1eYNzW4rNRKF
ZseGMG+th0lV7/+TM8JNSQYTnkC8qUCX4WB65FN+auYGzo2V5bWgEzDpsQ8GadVQcUlZe3I06wTu
SVjZ2NrJZ8v/iniObjyRdwrn+mPcop1/EDrPIW6O0hKhhs4jjXnqa0hF6vbKraszfgTg2YtgJKjq
1fBe1V4aVEEE9JVzYdKObgaiOGg3M8OFVGiXO2H5ML3im50EqVTv+fSwpEonxBFnrg+T18sk43Nm
WuzFwiAP5z11pbwT7Iv8HhEJl/f1exoMH5tjJQV+UYY2YF8w5yCcr10wON0L/JaUU5ra8oIf7YKF
oaE7rDSzYBjFtC91bJTKrZvGIqbkt0Nas/3qs7+p6nlRmem8AhksiK52AvnZA4OGxb1/0GsU07G3
JS9jKvGM3dd3Qiv802RgEMKudmvJcbeDU6zytlijQjrF3Dl1G2rtTwBXqdbluL/4fvqlDmHmgp1j
ZFX0+wBlyshUviduZx2OUsF19Gx56iqhlNGHC/8CMYnCZOLZVN5ELPWufdi46G3+NKu33HHk1XIe
vVMdkX6ZnMNgfVmrjsbx6XWo0GJlnClDvRvQS7c9bWOLdjEwgh63mmQutiyioXej5EcZ09wWJyw5
GVRNA6gdFkzhASMxp+LcR8jKA/28gnRZviXdSMQc4lUA4ldnzYvXih0NUW1vFaeoFBh30319whtY
Nn323DMlgs4pSkeMx7cq8SR4KhYtGm4u6SSbVEZ2RMcbGAjUWi3f153/D3EZcULWVrvKr124QMpY
otmS6urUTXLjrw/eCPD0ADHrTutI8eB/lgWSRxeEFqrTeXJi1E9v7D0Fv24b1kMEaMgBoT3A4zTV
eIwwsXGjhh10AGsCHO72PtpyBjpyr1aRQf64M9eAT4IKsnFisN/h2Ztv5VJGl612oYhRnynx6JaF
NezUbBJS7h0i1xHx5q/OgZnFxva0Od7hTItaU0lUl/Odniq+I8SxV3Gx++5tEG7Uz+Q002Pz/CWe
LGegohgL7lb9HVJETyjjB/QZD/S38MTT5eF7CBqSylBmNhffxN2Hvw8DHNbHUgcX/CXIZa28b3Vh
d8288iD2jSQeYpFBotBOXYbHOWSo/0moNxbAIoYLTgKJzjAJXDlq9fabUAnXaaTe5+9oUs+dwvJR
CzM6WMUkx7rRYN7Co9TWwSDwsrs1ZWsam21AxYS33pZcKhboPp7zNpsNZCkscZ1BMoflRnNI0MI7
JUqVISM8/aGcrKjpf7OVUbgs4DN0d7vo+W8M44M109CUY8A6MxPi/VWe2Ym4jbWJWv/yZAdq2fhh
dkuoE7iEsoR++1WiqGFwNwnsnCA6Ujhr2OZpia3ildnn2wBtSKNCxWMBt1LvzKbbUjZlMLqxrEvP
sqiiE9fantqkViMlIj8EtpxJBkRAuILm++IMq+vDriUDB+mNOQLNlCyubquBEW3yxmt1GpxHNTNU
J+rJ/AUlR37FXpZRbfGKUOvZHftUUSmZZsdfWU0/VlxeW9rjeFKSyuCwt25GAwGkIMyGDATyH6NY
mmLrnzu4SzUwbaep7V1esFvFtCpYRWGshiZ+BQHcCRS1VBrkAK8DiitENp6eKlvoVHn7XMZ5pgdK
u8RY47aaQnXcjyZALgzfGANl8M6pgxrm/ZmQKLnt2DJOJMD3dT2LX33DGKuiirSkPfg3XqNlKSiW
TeB7SW5rt1QuvKByWs85Yft4N0cD5IwZDNdhtNBdkP8c81q2Z9Qio3o/hRceUCD/7Qve4KohbQ6O
Qq0N2thsnq73naeet4OhqAcnVIiT8w4VtjtNrmRk348wSLBAnPS/PkH7J8A1ATfVkmbmBp2bJDNz
WWy8uCLIzqXNPDs6t92ayOMezKSTzzaCwK3Djl0JyIFtm26kT79RjkpdfMpT4iWkaERLx7nyh8Eu
1uHFqwtXdzhG7SFV5zNzFiKRREfQWBha7I5Pyj1vyVpYqTulT3b+GHmi/JBJ8FyPgXxdqj00n9xm
Tgqj8p+RmEWiqEhHwgJnABBejmWMaAsJBYvC1ABbdigpUnkqRVXu9ZGNzXpXpMgGRbrzMgX9VHzf
NCUMa26ZGfSy96TOqYo1TeBGqjaUz5TLMbhen/nuPCvvgyG/nw0nKQ8LZrt8v1poq6AA5WzeaEop
UIHhCgusL8iwEnB52/2JUXTwiV/7FVMbHdaStTS20En2q+EgnTq5SuGfskMLYn+DVG9a3d9tujG2
8FdYQK5cMAiiS7aMuSC1/vLRwB4aAtSW+YdR0aAy1u9oh4ELro8kmF63jDqsApuFpof9b6ifa821
0FBMFqDmPoDqnk2pOX50GEZZkV8tPAZU5J31RPjN8WVP+TRZl1j4HkwWt3dzArcUZP64u/6KyZ5q
rV4imDK11S9/ANDXV/1LZsSc8lr06cMP4K+J+iDhgBcw4bZ20lbIJXZlf6MEcfPzqn10nNVy7WzG
uXbROUcIBlUyJLj074l7vgVEdm7GeRdTSAMROziQ0pQig9+0U9/NMflOvapmCBj42ilLyqB7RB6N
WKvH2XbTGi8HVA0gBiEru5ESb/kcWPTIuM+4mSxtwtARF+U6X8PubsSnejEvukZvOkL1jMd6KpFm
9yU7WpQcR151pyi04jEfdEVRL8VO0pndhpG8VaSuX+VEPMLN6iBDa3T4MUOyswgE9XHM1wS/ZU8G
PEGErbxgRY1FSOOfcc7jqEq5OOOkGqMENn3OaaRJQSD9vK4JQpCsQMTJgSVUZXmTbUepoh+ikpCT
rxA8rBltTedEAl712JFa4WZ86lL/mZ4fbkuwSA3USr9RBufXseXziaUC4/YovWFt6OlRUOU9F+xd
T/77zrm4sPyTbWUE+bN3Ye+LlNxtF8+WLk3cw4lLQr6QQ6Um4gSlZhs1fpBxqZv81GbIPE0bykb8
peAY+WjbwOpqiN2asH3yBwho+09n8g/+s3lNMhJEcF5vx42qsvFBqGaK3FyxTNq2tCFYkOKNdGvf
xSP4Gv00ATBxOVT7hVq9rHUgwFYudSRglYTvU4YTv01g5z+djFbJicLBFEp4I8gyABH9tm7ChpkW
Rkf/TRJr4NBCr6kzYy/P52so511QjOWVMHCFF3PpJd763op4oIxVIruT94UP+PPkiJtjUIi8tqo3
arq37Wm972f14yezhc5fsEBPwtaq/1CesdhUsVPFXRK+ZOM+juQRbhksxeza/DQEVp9f8IOZjnOZ
yBi2GshUUf3el0TUATnW3oxrjNjYAbvciOFId5y9k0EbZlL9UNI8cjQ/XyfS/JctYQWKjWG/lsyq
0XWiKNwJ7GVgeBlJufyr16Fco+bE/isixM6pkFyD0wcO1otHHWrRyqx1OBvTwivT+aBqzOvwy1yN
ZhlpUjXzNmf4ItxgD9Tf8RCb3E9hfQxLzFaGzFumiCovwrX9ZSgMxMJR0hOX+44iK0VgPV0XauU9
GbGpqrqWUmArE+HGARc6MGU4jR4EgcUDtGregrcqyD1XE3Ke6/ZAUd2AA3BL7TtNncmMPBQvugQJ
mGDFN+yREN3rsujsPebtTtuLPbSg06nfkvmk4AsTYNF2ELtro6FrpKr1fFtqnCysEPbL/41beB0q
4B3qdvAh1kXRyGrGe5rBBrSwCpHR1FvMU43h/Qg1x61Qpu63BvqE4EV+U5KpkzYiiuhDteX+tNCY
hZT0ZtV+VqeG5XfRxUDHFOr5hZP9AzU0Nwpj4PyEvxdn2J7ijEhLOFga0QSb09Y3tc16N7QmxM9a
I34Lez7Xi32RUPHUo/4oCh6bpAlQI7smGjc7s1ccBgEp31eyIx+5lShp4YcgSXY1KG0cLEfpPP6R
axmOo4fsLahHRfuXSTFHHyz90xBwXuD6D2G1gattMjusPAzTzPyEUOVHTFK2VSkQiYu/uBucJoew
IFaE8ubPEa3AQ8NN9rvAxAaGkV7nPE+pm1QI5Vcxh4Iyta+Pca/s3EjKdySAPd0X7kTWhOVhDirF
hevH4NQieqChhe6zUo8hUNfbdc5aR3euq7ZWVL1TF/Gi6XREoM4AnD7WeAcFPuj+ZbwmMZP8GFDB
p8hxpb6s9w8sjfRVt+/urPUQlBQV3I4zhVsejy3DabbLx2PH/zeo8vx6GNgcNyaOnb7WtikajEeN
X3fDgQ3Fky9E9QRMvJd0aFdotl0SBQ0I1NktzSbIa2K37DhinU7pWbV70ve5GMPDPooMAdghsQjc
XBKFv3dOIXyWQRMaaiGYNGlSoSjCKrMQeevJRajqN0+xY0HoBLQkN4ioLbNvVjD8QOaN031FBaVT
3P1kF5LtHAdFNd2XYNWNytJ9DkfrMjqbV/nhCRTj5TjU80IZB+7/DEpOcBJNRZjo9bwh6upsFWf/
UeC9oc82MOo0/YtoFGZId86HoGL3QjThylqhx60vzKr9FPemEB5ZTnSJx+/CgxF5j9FJDMhP21a/
nHXoa3dpXLa1liV0b0WGi+6oABR+ygNg5FeNitwGk2mtBposVsLBOU63yK5LbDRR+jSs6HOv7K5H
sGLC0tz/5JBTWdQ6ue+Qxti5EzhNduO2NnvwmGqW0aOljPCKkEaT56ByjD9+TX/jrwXV0XAKgVHd
IpGNgBAL6ZBPrhOOUdk9V9/qNAazmnEAn3Eoo5MI+MfxkwjkQrfwq5fXfByEDeZ/8YrDk+E6nhQP
mzJ/LnDO1OGRJ3+vvmuntlS3CQCrX2RSvI+wEPCQl8EhHOodQYMrjmsKGZMBeQwRR732VvcOAe2i
v4y+gl+4TlyLYL+gJT0Cmy6k2ckJ7a1Fq3or11NqpH/0wejh2Dg3V2e+HQzPKl+eWk8dh8zc86Oi
wXeUeUj9VFbnJyiCsPLndNsw8ZuAM1qlzhcDrqCsPuJPtEUfqyPPNQnL4AtsJ1eEgO6s4gG9EI6V
h2pFAuevZPgG+Magur1MwF+1LOYjIXPdLX7OYSVqsrY5T/EISthvubMRXue66T1K2SFP83ZPOh/O
+HzzxdZ/28E9MAwDVCiwz50KuzwRjjseRmU8WGpTzt052LWrn9h7OM8tgRL21uWgZMIlDAD/Zz3c
92o0/KIIZWyua9NnvcjYA6isguLBTaA4k4bVBSIY6VLu3q84AgrIm+tgAOrjVQC0FRof0IWaKDpe
iSHa0yrvgEt6iYHViHeZUN3/K66Vd6hAHI8HzKfIdqT7aM5TlcnAK6M0rPF5aiGZ1WiCa/Yi6UMU
DCGPwDWil6ZGpN5ywuT9l92JZiXQyTAE0n5+ro76NLWBf32g1ZpgEhpkMGsTjnPgim9GQvA2FV2y
aZhOAKJruA1gW41ueCKr61N8TC4V27RBUIk4LpcW5KMue08ZTOaOEvw9WnTk7cm0nDFkWRlmRbBo
WONvQS7xfDxDko78rBhxby1uCr84wM6nXu6aRSJ8zD2y+rG62USNUiWvSrzYTHRjW3SucQk14f5Q
BiXE/HajOHMDFJsFc41ldw+lO/tqZ6tKY+T+LAX+MPc1ar9Z5OwjoMWbmzPh/jVs/5MMNlaUryBc
fccY9FjBHf19gu/6St/wYKLpdM3NzyeZ4rre5whf2713UpIHoXL3IlyKB3nQE1hL/Vm7I2qbU00z
ym57udb/MUaI+Azvdq29o51eua2jgZ5ugN+YB9OUVx9JiAv+WHuPWvQnXff/soqCv2OFHXfQ70wj
31mF5gavMxwvy8PULTaD0G1/glz+T1f2itRuBilaz8CcsbJqRFwHXKqhRcAbE/g+iwVnLl2nH0Tn
z2SzK5FdNZRdm1gCx+TzlULGxaJ01x2fRxli8x4B2568ksAu5PtsU4sMhh6OvpPMiFEjB5z1nCgl
Ddmk9PNdvlfMc2weu/a49Dsk8Tkrzyl5f8mHDFGvehOcfkrTrrhpVrldovyQw5p1+Xhhwc+LAhXW
uXsu+8wthWTX1lYf33Zqym6bJl2dgsIh4lKPRwXUw5rieq8kKjx+AKcmIuev35THkSSdVxhaAFvC
iQFRozI13am84uz2oG7fz9omtBVisnhHG/g3fRxbUm2ZojNosEIJlEKpaf2sngAO/kgmMwKWanXi
1lF14SVSit70Y2lBbUmjHPtuSn50Wrn7bNFfw/QDz3SF4btjGSdJ01OD9v/ZjLv9/UurGQX0iFQ+
6IGdhf5+/+mnKBlwNs1tWxEg36gQ1RvADLK+Ap6qLB1dZwvX4MP+8MBPQvtNV5nwE864wU2qisBO
Af1x/3qYNnPHFFNe43/ns861jtpdpCQqBd7ug9EjBDAkXi4K5AJK/CgMvEKdHMDtKV6S4nYlzZzP
QOOOVmf/y61N+x+v8fF7bHk2Jrkqqd+KYNUyXG83Dme7XhG2RZj8o6kES34wYj/mVDRmzF/NBy3O
lSaKJz7FhQ8rnYfOf8lsQpbBw5Hhdr78a32EaujOKpSY29InLimkcL06juEAa7uVL8Ey7RkeeLK6
OLliQJK9KPxdNCzfGLcZj5s0KGzIpgqX0Yrh9UI3Lr/eXk/LtLql2IJCecHnW/3JP5dII+HcjeE3
wKZaMflZRf0OVEowoajf37rkgwjlQ66yXRmh5n0lJSIMVK9m/Prou/uuWfTE8x5Px2/o/sre2QFD
9rpw+dGcWJeqp69FJRq/khnVfeyCG+ykDTMcr9YUHKf8XFdyIG6d4nu4EYjtjeOj86PsQnYOZpci
CkZI9J/MrxvOXVMb+IgO94AaFmbBhUDud+VI3CngKnRlj88GEclJA1wdWPGAFvDidgTHkHHOyRmF
8ve1y5LsYETFWp4wvshNQXlANFtyzMmtY/m45RcABrNIOcId7/f+cr+TeOJvRNw+uCBUDbzAeo1u
wktigpf8GaY4aWg78mXJOBXNavaXQN7IZZ1fy9ihEF0xtTSvEbUiC4EeWM/9pcJB+VPERTIuh/od
XRlZtlmWfKqKEYL/vnGPnC53HRqLHzOMJz/QwCLV+NU7+7UoHiD6mm20Ck6tROdny2YT7GO+GFQh
3tgZ9GWlw8qZBoS4JOuLAc2f9YWR81DSNK1YlKmsNoeDB+IHrU6nndP3FyUgJRooF2bmD3BuZIvE
dd/A/i9WB3baq2QxaBnmX6HmfbkRinopaC7drORVPNWmmwL0usqFCBRL85iepU/FHMUwrciApA77
s/Ji2Hh7r3NrBMzuETGdp7H4gr0T6nI5o5C4OIKJcNyJmwwCVQn8LObqpZVFjvIb6VCZRmY7+1Zg
WUm0UdBxXrESr1BocxarD4mVKUSEKO8BZxFBOzgZEUNxOdkWfRlweO4ufLzhveAp2wFLLK1zgY3p
5KE2FsHMaenlxYIvNUa5bmu4PuRR+gxK+Kff0om6njj5Fjd/FpbRceYWEftoWiHOkfaWyeBvpel9
iHHwvJ8sf+mUmITkVNKrUUsD2WNhcarA0GUYY5P0jtS9iaDt9H1fLA6aD0SNrrqK0jnUZtA/8ryA
b47EgJuzYdp6V58aw/3sTijYKnefolClnYQbxV/ch1G4HtxNEQDqCw6lRbNeURp9cuJvKr0fIOJR
ZNsJsj16qB2XkdQjzvkItR+jmxP2/5uJMIL4LDqb/oOWB5LrW5EgLdnOlQ6sC7ZVLD7XPeuGqz0t
30eUVa/wEp6+M1voJiBfAY08YaXFzK/Qldn6tx/N5mxOS4XIksw6zyRqc5L12nFm3sczll3Vc3Ju
WTb48VTnq2ft8uxd8Ls+2rFisElqXsIa6m182f/m6Krth9Mz1h8fXKtz+TUJR858FdF2DTZX3Klf
qvWnbSWts7eTzIMVcKqWDCBch52wV4W8vB6Rjr6Nn+9KM/WwGapewLTxf93AAL1ITnln49RZ5P+f
0/pd2yt0HR1AQHy6Iab6A09RIsJW+K3oeAqQbud9ZQbNmMVl04CM18zYWFPZjxW1KGPK2A1qhB0S
8+kt6+5CTTqZvIpQstlFsSjv0Li3celjNDFISkUQgjay9iMgu2kQfUxx8VNPvl7Pk+SHOLq3eKNW
WNpLKc0ZEUJLHs1r2zpNBVQxumZc4jBtwZzZrHgRm309kpdBUYhd6pWxV9wEpHYECztPS16e2dSC
BQD/WgsfLrND2v6Ag8GA3GuIoXJmHk0ZuoPYrLBsp2/KWIyGYeoNJxqi7UQB/MLSee91W7k7T8iK
81TEIleeEa0aTclOIviDRL1yKg+cqr7J5FQUX7sJl3gsH1w1DpLvFC4FoI/x9BRjFvq8ImPtqOQR
HMS8h3W3Zdh1dHjPJn1U2tPMH56VzAoHGp7K+DJNmJrGJa9HJ455JzBFnjomS41J9UNCwXn3EGB+
8Qg9m+itsBBTj9/ytXawHZF9xGmQjUnY3Ed+EK/cqcSvg7Yh7CYHpWUA8k/whnCB2haAX8xlwkLf
fGXn5hyNJcAt+K/4hC0dIlLdbUGiDQc6JV4+P5rQf1tXOkqxEUPz5usnc+WkSrjvYrbHRoCEY9iP
iu9NohstYuCQ6qtpRn3BJzxFYPDSMWEYjNkZkMiKvv90L5JqrNe1XwRwUyBnuYEAI3xjCWqqWzL6
jflPZpQTNEXcAJ7LLG911k8RI7blo1k3w81NsOb9ohGjR3jw3h7kkoDru2u0ek3TSclz9vF/3bU3
izU8mJxFEYWImyJpW9q+JsuoP3zd+U4Nk06rVtWDuWIau2NfU8M3B//DfaBHSdT4pBmqZrWzhLtu
bd6ROsY5k0PvuaEMrt7kU960Fzs28L2f63ZXQOGpTlZxRuAfJWZc5DXOOmArHejegbme93mmv4cu
l0vF+jXY3AheUAEN/HvN7uuf+SLGx7PBCii+rbfgFkQLXXn+O/IhSisKjG4XFFMjcBIDLDnH6Ivc
fHfI3FIBSzn2doQOusrdGa+qyAcTSMyjL8MUFN0ElBTGAMX0Pq179DjxS6Vrbm0P3Gq0j5lUW7nP
qN2jgB+/T87zCcT9FnsM+bqPsVan0J5lLDrVYiQ1UF3Yw5u055J7vjX9rSin+Z9vFjYdMxGZ+ydC
JCLvQ2JAewaXDwjPR4pX5RD5beFz3iUR3W6g3XZw+V0dOroM26fdaL7qIP8mKDajVZOILutcGrDD
dDOx7CuNa73xNJEUs0/YnaxXvEqHAEDHnarsRqgjgP+v+z6keJZRHnkrepbYFSfvVyl6OpWtslSB
KGowPf7H8GTPLQiUvLEVB+5977PYyGrvFbKOsuOSRhlu+bdmh4uVYRTHgbZbyOyurMw2cSI87w2a
pUhakwz/IgnwD/jrlE2eFMr+QmHKcdaWGJfsntwptFFOTBEzqQ7Ak5BMPgXzMhhIBcGnkHJCjAD6
4jrbF46ZIoWKMeJ2Mc0Tk6J3VBEMW5IIW3YZP1NaFClS0BJZHdnIX4JCCLUQVZU5Qs+cwK7ScqJE
gZl8yTrGRIXt3AugyD38HZvsYkTOTmKmami1g14d28MVgFoR3VwbKVaLxZSMVL2ODF94z9xLwwm4
PMu8EEV0mu+ewWA+t3wI/do3ptkHqulcySCVvqYpOqJajzYmJGjmgI0VelpHFWQkBf5vR76ZNfXF
YjI2fMXDJEiQZvUNr6oj05vLqUQOzima8JqB8DjJjLpukFjIoAIzBBPwO9FxDeHEekbMFeA2+yit
9CTIaKea4fx1MsWd10pvpKhKOE6bT6XWyeUhPcZviTDlnwyzoQh+JdfQ/z+aPABkXB7f3NI5g/nt
dbksAV0wN/rRIyhVoZ+I8+aDPzPZ61S+UQUpsKQcH8C8eGy4XeskS0OGArVN4ydnChBxYudtolR9
o06FFvCXrpyMpL+YvHsHYSsHuQ5ETK45WscFgPS1MNKmrQFsWmrdGaWG4Q7H7oy+VjPHdsRbiX+I
3XwrpQyln6JCIQPij/1q2Rf3igRQ/j3JY9Cs/eCr5g/123ppAgKcrN81eYe1X2X7Kfa3W5Yq60f7
0LTglZPhKsc1+peRRRKA/m9pSjSiL4gqsq4E7zYzDW9COeVtxfcy9i+oUqPsGmzqc+tVy1WaNgxb
js/Sm0B4GLOg8BiLuGeEKSsltwX9vw/5Wh0tzOVvMTOhFB9DSzafFGXRTcU9T6tHRi+j0gpDZl5h
8mWRzHVcN7f/eVORmLm5748NeKp0ONcOYq4xJZKlSNRMtbxyqu3M9CqGlXnlUPqiQe1IuqXaRGuQ
fWxLIgOrK+aRfsby34owGkCOw0yzbaoMcbv/F1/88K2DR/bME5DKO2HVVwpdvhk8NSHgroWy56WJ
jl/TOTCql08wXSlQD6QrZ2QlnGstSN2IReAJp/VLldM7AaIfL2CLCUD0CAL+WKgySxd87T9vghbF
yiI9fq9ZpP5eAXP99l7vfwR5D+cpGP7iclXBXsU9F1vMqPBuIfVBMEtYyrbQOTCC4wFFUJ8ckHOE
gw0OP3mFDCZRpjnG0c/KHC1YRcPmCAXMPoDK5zJKw7GnL9eWNpBpy++Zi//rmDuR5AxcADawP0+o
Kc8I8OKE4Ylz5QtBCHPnSDgdOCfmEeLQSbsyJCpFLBvGibwG/n4nG3AALZYzXprQkR87hWj9d3H1
KTtLosZ4vczLeJRFWRE1DrPdSBbPWaJHBPrvC0B4E3UxkeJxa6zkmYGJywRp0wnwuwvbsG8BNW6M
KsKJpd0FYddPjhAmRSKVpxxOsnkUjX4eTj0Evdc8GzL0be7UAjqZPTq3tbBFnMgQa2xiJWZrZBhE
4HeB54ziFEWCPc7xwVJA5NKr04PLEHf2Jk6Ae7KJZJgWBa862J26LyWwZKfF8UnyWG9qtQ8vL8YP
5DeED5P/MLZqbFUw86xZSn1Dgxw046sugSWcPga35a46BmhYxw1I15WOJ5DjU5JluY2dGM6yDruA
1V6RUz0aeMSi9RkhDgd5wu7FPW+bWLMgwaUlg1M3A37rFXZrYqiLDDBtgML3LBHQz1+DdN6g60Kx
cicnk4wbcrwOolday12Jtjdb7yRo5wBUa5FXvVqzmppvPDHZPEc0yKOxldlYmg/zYLUmOtSlQ0E7
24ZJccanm0E83wNkS3/GzmTn2RZlzDOuc8wFXKzIC2VBZhqHLLVk7gIjobJx+4s1KshHcV9DSFUc
uVJBt5GMZQ2F2ry/oajmUhZA+yvEdyAISTu+wEOOLYUHewOtXX69PrMWB4NuIm6CHxePhuyHfTJd
TUmitNRq2stctkNzvwCruEvGA5riN6O0btvgcWoOlsg+ngYqwhZXUCrFfyWgzY779NKgomu8ukLZ
lVC9q8H2Noli+QwSnodX/gy/XacGqYeDFxvJDqyPUXF+hKNE2MlfCoEFYOJj9u4Ug1xCwFXPpEt6
9WWC2ABO4edyN/wYYQGs+kK/JKbNQEr+5CfCmetcKuOtMAIMJASsoo7N/lz+8iAXA/tFVbOCqHg/
be4582y38ysD6UfMzRjGjsNNxg0+E2qLSsVTqaT7F98FP3+/aT7de699JLEdaKDwyj+Wb9VGIFIz
wftgBkZe8r5+W6UWijAQpNHtxZYo+Xhqzz9Bcxm5VtJu2wQmuYczqidOqshdiaxuDGKxZDv+CulS
zpS1ZkRGgVU5fKnXj0Ml3bYdserI0qEo5aOfEx+TVSkLnr5AuQXe8JwgPE/iNgucjRtEqIhyKldl
3mrchnoRzFTZe6VLuT/mcudDR0aIkwSn2TVLnZvhs7t4KAQw6X5ci1a6KovJLN85SKakAVG2yek3
O2zQyuP3OHIAb/nL9MHYiUTHK2Y0UlYaYCPLAwZPh5upBkQDaonbKAgwuZ9gO6vWBu/IbnZfLnEF
MiOs0/wo0pNob82w+CApPUEtKJBOV7pvXxo5jS6dexUuggG8zk8ZWI1kDmjmZRL1qZ7Q032wzpg0
UyX86DnURsG+kNydn9weDVj9HSknczxh6yIG1g4kwP1lPRv7qN1AfSmhUYjcf+hd3gg9Vw/ceHtx
QjMg4bbuQqQgyQCXb6iDkTzAiFdAery7mo5cj5GlRrS4uhlG4zg9KE15SuChAiXyDXetp50dnWgj
IZ+JGOVFapcVLLlSaCI9cxaAq+vGW+wl+Cu4dsir17A36+I5nziTS4qplWkYSsARTSyRWbcdPG52
xYYDgtlQow6eSjor65eW2LLbjZR/XyHlmMdRfLftAgOIgt2N+JOQVB3HnhA0jC/t/L/im+6hh+S0
PZDrb45TQywU5HSgh6t8JFBFK6ogo6I3vP3QbQyq19PZO8epuvyrOwu3RIEuGHl15kqajvyJMdZa
7YST6Cy3InS4a8EOCTZeTiYk2+1TxAPlbE/l18mQWoqDQq/vgVUC1Ex4kE2nxobc6QHC5ZID5UVF
fcvnvqnTCQ1qpwX7HQVHZFavb3ViyiToEKQ1b4zqHFYSiCC+cYTnKkFFNAAD8m+02OOzW1vgcCQj
vw4W/FPo8e6TDoysLlO4feAGxJlgENiK1VX/Hv0VJsVias29qcuJ6PAyRzRK85ISyjDZYem9/SOJ
4jqeIfOhKxIyO0El/s28M5y2jGnt4BeRMY4CpFXrjhVF3IxXlfEyFaXh+YGHDOdB20hnQHz/9qZa
xA6YoGXQBS68nz6hOPUrNvD7hxvyHpHyHSFVzTz/s2BpFvS0jjl0xMozhNN1oQZMUDZ/lPXibT5p
FoUJ29i45I5Vh93xN7V1h9ili62XavughJNgpnQTu6nP9woWUvbHCqGyKqrunifb8HRqMTBxC3Io
MD6RlgS1wwxpFV5Wrx5EA5/A5W+fhIGd0JLCwJt/ntqcfixzu71Ql08oyODTw23MGQqIjnTpKkZi
V1Aqn4ubdvm/JKAFe/RJEutNc1I9HEo5VX8TBNzz5eK2llfaSn/rygd/3v5pWoZlVuvOZKbpi2bb
6xxcnSA7iTGUHIT1h9doOrVf8yOFBrqIgMiFDQOs4EwmG88M+Nu75+tUPXN0SDOHYyrmL95Asmfi
AXOqX5Fs/IvM9C5FfFGLKISeyd6SdRC00zcwkgk7R9Bv37R5YncRbxZZ+iE3my/eltDkxtPG3mC/
J6+y3E58DeBasewt8Qldny5klLyRP1Oog4eFjKLY/XLGn+Uo9huUU87xGkrccN3dyg5Os0K2G4cT
6S/Gyhyrqe1MeaP21bkHFo7Z/UxVsUkaCNI9KmB4nuckmlVdOlzKVQ1jgd3ack48CIJ81d9JRMTX
1Px9ZMQ5p3we+Tg04fVfD7JMT0v3twvWshJzQoYMtHjjd6mH9nAAqqpuWIrwDb6C4688e3BjRCFA
nT5YRuSdcc284sQioflKdrQoGA3lOfRTq/dZ7W5D9Mpt50w1LSAsZHtyPHGi6YSLh1HyMLcYvw5k
FsvhQlFn76ro5RXSC6lX6C6kA77An8QXVOR7FSAfFBgv7coRvOA5eED/qXkeKlYPChdCXbERrIMr
vPKcn+dZhDcg+xFpXsGbbParAf4qRVzR/iBzSYGC/RyGdAeOtovcs6/Upy8HAzGp0uO8E6Mz2JqL
l3VFbz8gWaGRFn+SjEMSIQWksDfCOjlzUiV/nhBwTuxWkLibkJ84Xm171iB1kSku+DX5XS7ZUcfO
oOjleuBVnyXgKDZwk4ZCkg1KTfgsk+WbFmzIKQal1naGNw589giX8O3apqr1820ifkvSHIGHCHsA
qKdHLyY6UmqBlm/E1VHyogsbUtqTy2tz00uj9tsXwkDx7iBWARPKPkaQWjR7Dx3BCqCHT7Gsf6Hu
j3uU2PpM4fQR2EWKDg987BYl06Op7qv7uAz7JpJBbWsYqRWSGeoFwVQ/4JYm7XkoPeeZ3t0IITdP
3fAXJhc6+bstC5qcmIy9Ccsad+J83R/G2FugQE3OrncJmmE2AmvV/MgDJwVsv7J1f2+ejXdGR2tM
tSpdkvORhXHUzybOWiyYPh1/qxzeYeXUuR9Ey/OwOSoJaAsJIe5+w+a6tFlg265Mt5JlAQBx+79Y
R6f5fKtcLjYWzB02BMz9mj7fdWYE3CvKDtS30EQgf/F0yO5K3YHH9mbSz8FFAxAgeP/kl5J1s+jW
9nJv6HLhHJCiV+brlaa5BoahvEoY0YTR+MEzNamYaCrSEk9PsYz8LvT8s/q4Rust5OMn9Z3wzr36
VGNfIldIjwLzGa1smQXnj+d6kLSkgvLXbOWq7BWlXz+oUrKvAbNBwdqshOS44v2et49P4NqcRNsS
FeBMcZ2d5V+aiDxjvwzw42QiQQc6peB5bz6979eOByAQuNDNyvpP5kHi798qhY1BmL4tm27zF1vq
by5FdqddjOkPieLPQnYNzyiV4jbZ5bQXWZwVT0Om62XO/H3ewVIUgBpyeGEHrGZFfEytxsNGBvVV
VzsKeXX8C63gOqgU6NOEH4NHfzC5YIJYe89a3EIQ0Gd2eL3q+6mh3tqqPpXOB+ewJUDXybCJBsh+
Xl11A/ljveZIFUo2mS36bxgVKRcBlpIj+7ksp8EOAWswP/RQRvB9hDvmfl1Ycn1pODssAoeaN/uA
lU69bwumuJIjw3xL+d0H86TLAqdFxpXqzvJKrZHEp95FMJZMkvXwAIYMgUwe18TIZg5UIwkmmZe/
UQXH6VUELMKx2EmVe6B3BP5OAbXecCZ88eQbY2h4376Mof25T587tPF+0K4LLsOYiYv91K9aXTlK
4kJdy4Bt5rP4OvlWYSglSfN5P2dJg8iUnLVU/k/AZLotly9njs7vB/F4+XDg1ipZmC7+voQidINk
QM4Hu0Z1owAjRQcOot5iT2TeQpLEtcuRbgSaCLcN74dP15MpPtrmotk37PS/nxrR2Bbc3hARDYGt
5NsRg/0EDZ9EEERGQkBnFkRPEy5lTiLpmyDN54dnAE28r7u+zTNh/kgFI70dKRho54SVe3eJMZUI
nPPGsTVzCYdFOfX3DRwUrEezxXBNGnD7QWO1Xc4MZU1RpX529gkil98CfLbgc/Hf3iBewsUAhwNB
QYIh8wQC5mV5XUigeKo63Btoa+8VBL5LLrI2tBX2tDyjH6sJaPUKLyE0jmpewYG6llEUq0Lrifhg
rNYJ+2pgyW5VeaF72YhqUYoqp6A6mCbaVXQGL/y9XXTKw8iqh+MIag9eYEOBjGgevy2MKZK9zZIX
KXYhVKEl7hzjsucrK6xpW1v2nO4rABn1C/oc86E7UgdDids5PAyIq9yVFb4CGcX8EPmX/swaKUI9
z1eBsHp+C3pXCx3lCCb7xJA3EgtuT7/YSKg1U/IEYMMAEDTxHqF1aSEUEW9uPyvF+3MaUD3Fs7JV
MUnzsxdnmY/gnH1XfWIILSgrp5yUub4GY4gycCh8n1X4t2x7mxIRVz2GlMIv9R+81MkURGA8uvHl
xkaUS2vQaipcLm4xfdqAxAVAyVoWdlmKFYmjcUudK+LDrzoaZezgbJtcW1C16EYZJkRk6mrcFS+H
w0JA7D5eD5E1WiwEvXA/mvHb04I15CBDbgjT47TcrbjMSx1cjSFr1czaokABrHbuMCOYRojHHiU9
hDgoBvVOvveMBxTDx7wBJiEWZaWrPJe5aUi91x7ATnGhowmegV3Kadz2gIdx+ii4t4lrY0ojxFob
JaCKXM5O+fbpDys8q7mMlYi7pxq2cxoiehw92B0iNnSH62KTOUHprrx/s3bjZhXzdRP6uZSCUlN9
eFOsp932GOvkI70Ftjc8Dxh2UH4DrhvEEg9Y/i0XAEyu4mSDrwM9M5es44cHrTa3MfLPq2T3+x/S
GOhc4sf7FiiasMZdJI2yC0uYPDGUdpjdsYwqUx2Igxd0jWZjYC+rXjXPtHz8fNdB1uOSPFWLeNem
i+WnrcPx+qh3JG74Y2zeubrhW48GkLBysByC1MFJ7pwKSmmy99Tza+IJEsGbiVBGs+haSmF+roC6
lrKqNRh6F6BqhKm2TUlBuEN6+KvyrQFGL8ulGfzeyvz5fTNhneu+ux8rSyR8eZ8s7S+jZB0XBj6G
n54CI951tHz3Z8hQIW3scyVw3837q0xg7UflbyXNsFAEOu2Q8eONXGjKbjr9sBY8q9CYuqNMYfbJ
gfoVfTMUuyPD3cfXvvECbH4EGYyqk783Ajbyb+nP2j9gi2vSH97hbuZi9W3P/SeirJphqVI6wPcD
yVmcaCOQt8UGCtPmJkBcNF5dcdlmiwrklbEgfi8MZbQBWf12y87g08rF+o6+xqqyWBhLpLi0OLke
VM8Y19dpNdB8rJ9Q18PhC/wv8nnh2dxSJP7Kr9Xq1Rano7ye1g46URh1cIU2sPrH6oBJuRlvpBrv
48Ue7eOBheHxlb11SXH3fSqFpgu9X2p7um/T3xnKDcAqj8ZP+cuVTUCWJwC+k1Z/v+QGBax/fa0s
NBW51DsZIHBKboy25sXbC70+/4s7MRuVMzr6Ykys8Ohf5XgykdSqulLDdRCmoHLGyNWfCou9475f
B9t2Eddd5gsVR9boaOeQuTcr4fZOI+2oxRm4AkKq7N6XqsfaF+zOx9OyH0DldASGT0vMr9u2vlIB
8nnul+/bsaWVk/HsOSlUWPjZmzGQzCgLCts5ZxN6NZSszJVHHYYj708eq9LhE5jDG2Im3aQfi1aY
t/NaVMQfVZMMu54Y62PQSwHEp0unBKcHDrl65Tmdfcw9t7mhmANtcNXAyxcYoideQG1TEFnA8V6L
XIeSjwMCEC/aMI1p+4LKUj+48Us72+tqf9oxNNuoIWI1uz5EwOeKsIrKrB8Yx3BKXeppmlI6HVxn
ujM45vKqLO6Gn+b2zztPLUGMdN4cev+sGdRBPIJvCwd9IyekgpmLU1tSw7+lEZE3eirpgbIz6CGx
mQfr3nWqQhWYaH4erEQjDV3PWRyG8Il2/HGPL/jgyHxpgIGBSx/fdTbQhtSrBLX2VSDoMo/j027K
Hm8/TgGQfLnT/T7wj6tOhLLLEgq3i6//i+wyU3cIUdV3a5DtlCsZiy0BHGzYJoKmcgVhroh+MBEl
ev/42kKZCTFRQem8Zo75pLl1vmD9G03TH9r1wJ7hcDBtX/YxjWI/niFajItXxj6Pxkriii7xGHKS
Krz0KCKzCyEJWgyFpDsFzygycwsIDfZyJKspl64v/g4b2LqU+IcVypvw15y6ycnw33vZlpJU0Vxq
P1etciMT41VIVMEr9iBGS8g0wNhiN2bA/rOd+DH+INF3fo4TVi3Api2CDIisPjW14JUu3Rxs4KGs
lIRaFNy+n493NkadsUtWidJOEepRQWlFGM2jxVC0hT/UBK1IpAnPEE670rnLZlN8zfjBILF8NFd7
MprW9ELjLgFisjNoeF8QnW8LOSOiHcMDM9ze430WR9KIxw+h2jDoaFq72YBuhd6ZO/A50jpgRReW
fehalMM6ZSarKO6Vj7yAoZG9vfnuT8yBDAW1ofYGpyPcbPRJmCUdDCQNBN//R8m5kM0da/zgBiV0
XlhmzUuA6JLgsmz3kGneNAUCJ10UENyWp6IKrCMJE6MURabnLlBILrX+1tCLD81Um7snBiZQkRlk
jG3UK+rZtMjd2YmUXCaaQM9JFXWFRi+AsYysDPBr+dxJSVNOw6T5f5MixtsF2NnA3JdTVwoMTOIe
/uDlRmC86ZEgYQt2y6yrtb7fX2XkT2hWcH1pZj9WHlHGmAM5K/uIChqgoJjXqbTdB/v0M0b3gGsk
1oJGaAbo9Twn7zWzne8bVcnZkjtWlgc1/U0VkO+C110fNk4HUawuC/Gg6/xWB6Nq4w5eyEmO1eT8
BUGkYNajIxkUtSEnlVXBm/WSTYZOZpAP1bxTSrU7WL5sGwBZmmctN/Luh4toZ2aSLAE+sYu2bLi1
0WuvgZMETobShnkbkL2Oniel+9YufQ4nrdofmss67Pck6+MKE5SAyjHlfdIDruuEzPc7hbUlipbg
cTDBxi1+ihQp1DjG99c8smrIqWWrC4RyHrUZZvUcJlieWH6CoUnlYnOO7A23OGMWqSRnKCptceHd
ZEPAi/Mj2Njgn5sLVDBgmc3hjnszZPJ2/LX/VJZ1ks3ie3O2qK1fZwaxjnN3+RdbYR5abIpHleJ/
MSwPswXLgPhwJFY6S9jjKn70PztcqGXpQLU0O703ML+lLFlLPntHQwLraoczjOLguZA7LM3k1KVo
KDAlrv8RZUNrKgLSVevto7DjMKSvxwdfEzt7vfXtuKZDMK5bUD164heQ1GVTchB3ygOLbiEam36l
alLS1DcoaM7mgUiTMNEH0qa6v3zA9LwhXEMFyFGw0qtbsFdV4ic+MKpsFSqgTPidfgeaHNw1lho/
3oW7U02wb2EQWZ67cDmLBCqumgV7Q6lX6t63rW9JL1qIs57F7KL2w4z6jUVQhgHBjDTmuJ5fYotk
yXWqrspYtUWYj2tjaSOu3LC9R8RDKQ4+WRTchbSQs0e654fFYVp07CoGHCAlnWPsPsTYSm3B3PNf
C3X4dHKrLvCo2KW+vJc77LfvxwOFxLIC0Fdz7zMrFB7icJIr2bwkk8Zkf8Xr+0/Y2tsx9NXas3ls
vQ8aByOcfsPAAl0oZ03iDtQ+yxP39LWnvVpHpNlnE8u65qdyhzOlIDg2bflW8RwP4LsBfAvBRCFf
hA4gF/c9jxjyovQcflE7jy1DbEVLLoQ8tzrNvv6uPNmLoy6xyZLMwiXJMj1dbLd6o+ylDqcrgJUQ
clOlKlKD4zxvsjJokDhR6kLp4yH9+Y8TQh+Py6LyaQWRGONynUljxhiwEj0z1YddcgFMW1AGyeFp
21fZdCU2Fe0tSLTH79+jyZkRQ0Z2oPhWt4Idb7NQdOWfG6bMu2rpstYmiH9WKDOYhSfm7K0VzaZy
sHAGjtsK0d0VKhZ4xFDIYusoe60xhH24VR/3Fjb+sxYD8AOWehfmKmi4S6MBkGFLw50zBLvRcYCa
AQcQY6nA6NIzNif2p/tmidMzaU3t5WQ6Q3c6iJH3bH4TNGUz2uRpuUCNNzvZK/iIqNkRikp6GDUh
VnlvNbgE3ImRrD+227TSrPIIOUvGeCXX5R+U1j0a0SYEafo8WiUsMbU1eEUUhW4vq/XhAIT8Vhkd
Hv6lqiFO+QchAb1N5nsOG13q0hnBW+16P7ZMLkXkUeo77ZbwlOdzsmnTrhb86ux0/oXzIrqRD9Fj
aIHZuzuRTq7buG3XheuejX1p7DOGH6IcJJ2UndtMjk62flkJdpDp9sS5r3I2sKjyq2RmNOzW6tD8
Y+Ec8RoROLXj26F+XwhyTO0mUjtof9W79VnWSfLzDZzBatYI4JOcmUgQjgf0/V1udosFryrhJcM0
UXNssXdqRqY8Qth0wiPokZCIyStMDvDBG9Na3XcepGv8V+UUlznfHrGOdqjUKiWsytPVFIOwYwE0
/QKouyVERizWPQTSTHKQyhOj2zGYP9kNwQhlbYtH3NGZ+iqoWfZMf3n5HDVrs0asohmVJJ9qmhy0
jwGlQ4nv+PJ7CVFEmRkaD1d2SYPQwR5uO/lj45Dbzgav+N5Sdm7SOUWFXLLa7b5NqwoMeNkkethB
2/d4MpeTmJI5XjRdkFb2IMjuQZrrTfatu+PcKZM6g9EKRBzfZKd0Po/8LHWYbqQrq62FJXMuXpob
5RBMlxyJiJ/K/KYuTz1Ht1FmrTLQy5udZJTsi7len47wdMvNqTs+ngzfcWIfolEeh5JM5RlQNN69
oxPHYrmHnOqeW840TWOoBIoLwIqngQxinNDArJzX7kgTQhFZoNzMw7eerC7s8hP6pTbzH9CP8Tzv
8XTXo9k90k7Fko5E1fTP1XrnOJKyJuEBX1f/lYJjleie50OzRNDOS7XOUj05T7OuFHbbYF4QY7TZ
BMYGyGzpFNFfDwNXFxWda+tcaYKWrY22mHj4o1CPO6flNKtOwmEPiNKi4Iv9tFH7uialqBT8tOSr
HSB/uTA0E/z33pMNV5PsiV2k8gCE2tPOwV/KxiNTq5Acz0XxgHycBF+6Wl8IpKw5bJ5udWwLY/+i
KzuGAC5LJVTvLf5CjbdrEhIiyvAvbDenemKxj0Wj2fOtQkMA9MLNp7Mq36Im+EKm3+lGLEwbujVM
6+9bQUepyubZ0yCeU+PZOjRlQaovxhZI3l7aAPaCIsEBsTtd4kKfERIZOwNvNqZg/Yl5IZv61k+r
DmsIuGkdzAJ6IzHcfPFzJAI6LmcVwJiKDvI73xjgvvHRMZO9O0FIVSGLbBZqc+3v48UgSM1qjurd
0/l5CX7yli49mZjy+8XXL9RHaVvhHkRlKGQN6KI3T6a4IpXlBZtxZLLXPzsl8rZ5A+5fMzVCEaxe
MxybDuk3Gd15Yy5CPtuC0e7sLrpBuPKb6V/zktMPwBbXcq2EChJCH75P9sgdENBWodb/SqzIwc72
PJ75v6uWxtRr4P7UH4AoxJKUkWcVCCGf8rvFpq6Ts/+e7TOKIT9CrCKy9NVfhBvmqAaJyFCTsf/M
e6xJ58f6kcAL4fASjDJzwNcm7xdZ0CDj5SW1kvU7z3MQMTxnh4QgsMM62hL0gzRue4NQC8YhZtcY
BmO80Fqwq+Mbm4tqd44m43C9W2CzPWoIvN/x6JwcI6FPZdJdHzPMurqsGPDisbUrAAYssbxLjjQx
88ri/AYTd9+tzjwCcbv97iG+maZ4ydYympgZUipmBkJ4ArTXf4ty874bczt2H0W81Oesdd/bN8j/
51VuseJn6LYrULC30fMF8TRG7k06/dWl6GF4oeg6sXcbgDIEH9JYpIWBk5nOSjh6iHLiRxUyr8vW
v6fkZ+pHtEA2tKOsrDXsShxefm/eFYn79nqtF7m4qeVMJQ2uxXwGFq+SwL7xNwVRXbJpecEFQ5Ix
mNa7XoCoMXCaEGeCiTUHWKVmFsRuptw+nwh+eszGMEm9VQ39/wNCsVWTO4NxDwnDbId0yU4Se5BZ
WZnxlmmEnSsd7lyTUEXtWUVyFqYXagXbco3HlUKEMtl9fa/8w8qP9gXEBA2oi5AjUER0Xc++AbEo
cIRBu0maf6dyABaX6ZPJq7OdlIjMJZEHS71teBs4bLS2yXxDtu9/DZkFpFQhGZKN/vuKI/fMhj1c
2pgZOwWdkW9R2GsMFg+cHoee+aMnodUF2y2h+id9DRA3TK8NkxIzMBTsXHFJChL04S1nPMxoVViK
2/5bJ6ObICc9eLL5F4re/Lbz63D/dzjaasKL3b1RvVA+Xpna3QBTV1dEgk3t1vjdvC3zMqsJAoWq
SaXJESrSF/A3vSA4xBQl1uNB+sXohMylPJ4Ek2ve4qm0SVaHv1nFmmeaV2zhNzNkaTDushVZl+yo
zZHqQxAIyB8Z4mUxw2ul/insCN3SDbrhPJhHw+pIj5KW+gGvxQhsblCcG3mzaJVJpj0/qezx9NNc
KMVZ2Lu3faGyg8tI3LzslbS8+7QgWjOIeTUCcXiwIGG2AviBIOWBT496k66ktMq5QnmNs9KdpaoE
/axjAg8lgbk+Hh/08nMzT0QLAyvUY3Frj1gAtKOXNTx4Xxbu1R7YSE9Iin++dd1X9PQPA0I3CUlv
1xbO6WFQWo7x+n2VEPA88uaHgPD+WkQMSR7pCg5gGavYSEmpXcpODYMAz2isf//s4TMjnYvOCnMJ
aVHaHsFXGgLNC+6pjkpTQR+lUDHpI559Pf8q9lryHJPXtInMBEjgzIpx1bL1MTK9XM1HgEy6CkIU
2ZPMYhAKWhL2xY/Nrhg/QldV1xkdMrPutCluXf5wcn3BvyGoic3bNwl1q4ZGToc3n/ypgulRQV7G
5+oe7qT8+JPSvT2sgzn5Y7sg+/A+ToXC+7gKWRx+ZeaG0rc5yGDTNqbgRsFlkHKTVQ2IDFOS1Yrh
kNJH4XeAPWBVP63Yp+aMMMNXZRlExzA4f89NWbgyPnVpmvf7PjLZDGZ3qLWeWKtW6bpss7Ng9UKV
7ZIAzH8MRkocKrnCJ5nl8fD4r105gn9Pq3Hq2ZAai0fRfL3vlFshzMpf24UVIdL2QmBxuxgyjuE4
ATpsVLw6ckS5B+vKgHVhArFlw0VurRQsTlbdOry5EyIvs4kKnbHxn1e4XqFopQRSRNhtfwV+TLiQ
jp+mqLmSyLIGtyR83X7j/sRKk6hu7OKtRTAqIWmWdVg00/2D1+GHvVc/GpObo48LAA+scQ06qK/R
IGYGW5pZ0uRVAilLv8E0T31MkkdMyu6/rr6ANcvQLokDA0NQpN1UfyTqitKdkF8+Qil9HiY5Imbn
p1tCOeatNtZ7+GVKgy/eVyygSUS+M/OsDP1pyOax9czJ8sm5OU8zexDt2BmAT9yHZ1NbCTCljZTi
pZsyIl0o/Me4+Y48Q6+KOBYjEXxmlAnoZTgVa14fDi8tYtVa/OgfximzQxNqmtsmdmovIpn+bZIH
vgPGCqBfqaDNQc1VPOomLHFn48Mb3Bic3/SSKuIhLbn9hc/VZA2G8fzHZabqbLH2FsM+SpGW8EdC
ASVg9po+1/Xk4ZGiFly0Ms2ZPau6/G0Kv0YjHfjyU9HDlraMjnLcny1CqQzTAGxmiRncJI7HYc29
jY2eZX8fohY5U11AAVnXQyM5Uio/6CsRsAoydqF/FXVcV+sHCvnGej54JsaIebAHb7unu8MxzTw9
ppBGdnkzsYHOF+3YYCC7y5mMBe6XIxJdpvuDjmz6vFByedAIQ8HBo34CzSjpI7/ivPWduyWEDmE1
/i7RPFVHRP7SHhVx1rwfjMBJUN5vwwZGjP1ZnZKDVZSiiiCYnwM3fUITmJeBTzWpOG3BoPilNMre
2n4CZ1+yt8Vclgjbf8WweiVKaP8WAwP+WEG3FgJr0ZZFhNX4JKTwA8u9/WxyKWgDqNewHmrSAEaJ
qMiW3sPUDFz3XfVROx+kxoLaBvTEY4U3QeLzpJMeHteZTZ49SqC+B0ltyLHV5W6Ee5KtSRymxIGz
EqwV0OOtdSA0AQG4DOSA2afh//dvVNZRziqI5kCbXPjTTKZwHc/1iFPl1Rcdgoz4kTqSe7HZtU3z
9WBkHeHJKXB7mnAkTs3j4Aaz4igrIeI/AOrV7Mo9ZK+mZD5NSjZ1B86pOJkh0ssiTK6mcvlyxUFg
if6eCAlR9JjsDpznej6NFkOe7Zf+5Z4w4q/rH15gNMV5pySSTritpkisn6kKNjoiC9tN8gFodoXp
XTWcHtZ7ekrpfcRR5NSvLswDCdNnLG1+VcTsx80Wu90NQ+vNkuhmKPP2summOMJQe0+2QazBpy08
sxiqp01DlMgQMomtFicFmIl80WrnQESCPNvRS4oU/WGeOTMAARUGv22TUTggxXhC5lcpdGPQyOQG
csF3NvcGV4HL6IP+kgionylx/5OaMvh3xbhSzvTRkeTiUhkrkMWDsp6SxaXYA4jQh9pAdh1nZEls
Z77xD6QbeFB1gKV0rq4Oc3VZ0JG4Zi4/kDF58+3Ysk3wCGHEB1TVAmh+XFMzMoW11Jpx42zB3lFW
UhIqQcXq69Zx59SJjjtVdVKYPlxgPxQwrf4YyVWJ9hB4WndcG0WWVplVPYuuROfHkKdCct5e69F1
JTH/1n9n0z5Efxrv75CQDwOgJEm/QiSzH3vm0x7Ag8OeKA4slUfZCjOFewy3gTcbA6stCzwwBfZG
EcyLpNggg/3o/hRFxVOe1DBR2ry67BIXMurLVwiKbiNCnAml2+msPUogplIdKGnPGiWQU4WO2tys
Pb6Kq0LrIFtdzDtkIaSYBfaIOHGLuyLD80vUDG8rPQJmE/UKtZXxbixA+Palme7Uyzn7UFuO55Cb
6KsRnEY9ZcY8nsKWKc7fhU3wPQkTXh9jws3/tOSWjWDa6iyeQTuo/PnkbE5CebJCZ6tGg0SGF+gW
J1qL6dEQHbMpXksyMy3ui9it073UKbqFDQb6Zh4yI5gjlpLdKT/SEAqzOopTsnpi5aWmwW0AzG6Q
//y6VUStJ1rHwCzaWIIfl8E5WxrOi+uYZ994X/1PfeeW/kjqd3PPmzD5yHAuAsklyha8vQr/D3j3
sS/yxodXnh6n5ZtoiNRxrnUk/07WMQ1vfF7mVFgmVoVOUmAGAZLO5VgO1+IETEm5G3UkLMmtr04t
ouWc9Jlj0Dupb00ZbK5f5W/ht7itzUqju08leHw6Se3X/7M5xMFY/l2WEBPNHmh4KUtekv99GjBP
ef4Lq+xV1ki/7AgCB0u69NNwjKuNT+FUXW/snsmNe7GD/3Wq1brjt8QmLbcczObguhXtrslpa+fo
IAB9L4axbRXoSRO+/QXlpHKDEcUSl5vHFyLLrQqeU9Xtcu3B1bcKL/tkCV9JfJWwSOZdge3jea5B
Y/mzVIkarXobGq5PaUNeg0YXzPo6X7l3WCFWjZtoZri4BnTF9/cX/dJd+q1RjOPkE9GapzmkYz6o
rvt1ZSydW6t/T4gSAxD7PLMbqkS9kureA8zVbVDkUdDhJmh4KDfAuU3qdOq/JZKtfBFGTFJLgSsT
3D3BUaf0wTipR3AW6zZFhQQ1tDWhLBA3imrkqA6jwkT5xmV2iGbvZoOA9IJH502WV1zQZY97wewk
P6srQuDiuze5shA8XpQ/F1Jz2Ey/rWB5UJ7LgFsLGwWVzTJUBPO9TRs0ePHoZUh/LCwn6xD/WMxB
PGDLLfVuT92uKWPZmr22lYc2hifNl+vqyI0oKbKraKSl6ioxNdNWSlOd/aAX7oCvC7iJB759uaHx
CVbkkYudKflaxRlLRfs/1oAkjo27uSsJTkMhObuIAPf6o3IMBBodyphFWi4UshhmM61a0US6yDbt
ojXWYjZcWlunRXkZLTSP3ZXsAHmd2wNG0vBkno7Qah9DVpyo3IeICcjP1uAOVafcDVOYP4AsyX7N
qLDRT01Zw/6es0+x5CadTB1i7nf8uz8fj9GIXvQc7efB/8R+VJXxF7UXw337Yv5814DYm0Mvv98W
KGFbGhBKXNvsh7RY83VivwxxSjCafEwrtByjNNSxtzOOncvmYEa0vRWDfZrGrB9NznAK1+c4Nt37
p7k6Q2tWX+PQdqFj5WJ5W7tm45mZaGYlr2ywSMPtyc1CDmY/2HIEDUHHBLA4Rx0/diwwxl0bDu1+
ySUDgrI2x/ZmRMdw6hYvMKQ4ohE7zFO3MwDRfdcsv4K2/pTVmRD3ZB/KTM2DqbTg+yieq+et4R6e
h9VtH2Ivcnk7cQyKqk/epou4abJXBytH6UMdRn5hjki9N60bFiZdHicB4/wt9JTYsg8EuB+fjVH2
Cb5QW6BCROI/qKghD6UGD3jSUOlO48avptGq8H5dl2JnUfsxvlInGsAhkyyml8e/Zozu7cLgepzo
Sm1dFWJSGovzlF61uhvZFtIBk7GzAtO1ecwvw/MAU2R4X82+iisB9oZjYQ1Hd27Mgpx5QQoNYEd7
x7OyWAliPODbV7DVHlgN884JjQisUZF+yr1thXKVs6BrEZSPvYYR3g4F04dMTaRr85358wAfN3Cr
2NTZ8qnSFiO/A9C4IMHciJp5zOMRe5d/f4uikyx7E/kIknGNnxCV/7PedMxh+U2bkyMsXiOEv9yQ
6KfjKkUALpAvYNxkINzeRAPrYXwlyV3lPR1IiQ+CQZ8FOQpCcLYrsTHESuRw6hT6E8783Afc/gPR
NLU8HnpYSttthmKLsb4DMXlYVabNv9oPMaSbpQpQ52Aa1srE14GN9GwBvU+5jKJPx2qvs1u0nqzx
93ihmufU0PAKB17pz7SqzGAspUhtpcjoSUQXqyowF6kOKfcHQKUq/zJkkzm1VaIPm59bdCZfnBgw
Z7EbFnACCboM9mr1gYVAC25Ykt0wHeSKeBIDVKd1NOVo6rL8W+LY/IKTC13+1sL+iXyh2Ev+oar+
Zsb/3d8jT5MCM1/BhQOfG0Nv0EM0Q6Iyo5v6uDQh3AfOCsx6SuFnZ9TGumYgSBYRojdkl/Uzk3tm
UvtvabPboPQw5UhDxpGnjyraBnJysUH8n2HbREVI7hBkGbrB37qTwJ1HKDvN2n1hhOp0Kk2rSDH7
QIPjagIclFrHr3UuxzgGSPCCfWtsS+3GsC58tuDUqet8JHULsBorWQE3FTq5nKa+jS0YCjKNSlie
ceLR00Df/VfZA3qG+e4bYUBn0KKkmDQGdkfPevIye6rB8gFZQROyQ6+NEYBKUY56gEj5H3GUh9cQ
vsvtiZ5nJZBpT/rCJd2+RITmPb874EEaB9XSD7+AhvMrJY4YoPD9fI37DVpspmbghECIncKW4Bm7
Et9Z/g7m7gchAVFx0qER+p7j9RhSw7CAyVT3xzLzvfft7sdIdgVUmhRfiT7gc9D+CY6DloMAHOi8
WVHWAFTLNAqQhfFlg6gtMy8p6wgMk2hstTHLklSgU7T6g1v6Di7JCYujCCLst6xa1AErtaz2/Mw7
ybsMOFRlI4zMYLnneuyEYGIPU7U8uLBKwodkTwTondeDhTniO7JscN21+oMYRsK5R8DuvZIKjvJ3
NvbUeI4BNV4NRbc/ozTM9sqNBgIa7GWxanZovR0JAMqNzVRS5cThg+zvUb8AUrDuQkuRNPdfXqWz
0hy2O5vqkzLs5BvPcKnc6wVxrjGesxQWK4rxsir5YFYE8HWdz/ZkBZfGUmnHFbXWHr+R3Us8FBun
lTKF4FGN4UKQ83vjPNEU7BP3hAW3+XsoJzXXlgLWSB7UbrpAfsfZ1C5IVfpBRNJNSmzpBAMUdhMw
m+XHEAC+ceUGkElaVcd7PRpvuEw1AlAY6uDNY1drWPX5BWPlW/1aqAt90lpfhhBS0XIoshwG6Tyo
AVrWnZ8XxJHRbMqfHBSmE3Mwv9oI2KwESJ5mstCqfM+R8WPVKa9MD6V4ydw8G5aOccRCh4kn+BFn
E3TqKLNUMLCkRBHJwJUqv3gaxMlHG1tXz143ROzMmAKI67SvmhJbxcIrhee4keBj1a0rtaU6jX9p
f7xw24h+TVK9+5WQv7d367trgUqAQnOEnL8SY9dn1SMmjzXKRJnNzES4EG598pA2ZPtgz9Ey4l+X
fandJuF4zkQ0PZ26dRGa8Jie/wDXWm/lR3LAL9ZW9dsiXNRJf8t0P8NRoVqX8TfBJUvTUcvSQLHr
ZU+WjF67ijMoHXRITrnmbAEuERBVwwXGSUeHntapsMkaxrM9PLzsmFsFAByhL20ZchVfS79SfoXE
OIhas0c2668odixY2oORGDaqF7rhaObdctbO26/Pfywjnb/wZBIpjQXRnHzglPM9SYN9mfS+6LCk
VieHCGZcn6bANrAXGMSw9oEVtX5cPwTq+f/8VBDP3v1U8ghzZ+WqBnfcg8jdvIfgVgZceRiVDjWE
qC+QpKPHgS2tFyN9kGPcIe3toLl/GaCpEiebG6xhHXux7pAV28oQRXfWiWq3RG+3Hbh//+P/a3vR
MEKmX5VjB9duCmzmo+7HCCJhlRx56txwoBCfqQ/85midwreGh55Njf4T/upfmW7+uZ0WXnuCNExW
22zZYizkUJfjmj15gkDmN864VzPHiQAYyWcvuEt+9c2n+Xxjx+BwqYw3X88wnXlc4p8jui2hE50C
YI9CmExBuEkMoO2wCQxNWAOjB1MZBWbCJwnkP0gjhOxpCmqQhsTkFQgU+F06LE8EB3m/G+J4TPSX
SyWD06iAJuZsgfJnDVUQcp6huHjfvuPvKJPY6j0B2IZrzqo4tpHQZikcMCYUsXAleWWPLuIoWXTY
2us+L6+6ZXAd2CjoriCqJyQ2MIU3TJaGMZtazVW943ewO7p0H46uMIUE/u71B51g6ncG9+e/sJcR
JZq2ld/SZuRG48qfXykdBHgQYY4evMEs6VTjxqwGbRTj7LOoiEo9gYXle0trApjbQKIlBsYRp1Ib
gGWnwgP1OI/+04KhLGVjR9Fc8K9ZzVjJarEGD/TGa9/ozSkajPviUYlkEAKonvhhRfExz/LHVSym
0YL5VSLaEC4vJ/zO2PnIpRAbrMgyVZzKiH89HMBsahJLuSfC+zpBZ7HBLOUZOQQ8u6PXZrkPtLWr
HLKzb/OELhCeZMxZfzk9cHChzjhlwC0nb162JU/czZUoAzaKZdmL7UnJPBH4JAuDQWKNeNvkSdHH
UZwwwjSdEGNjHQITQ9+VEWjcjhtkX9QeW4kqEpEqkJTnOpwb7238dIvkENGBcbpUBXurZgAyr6sA
ImQNUMTYdGGrPAZ5nvMvUEfiU+tmRK7aLeQXKGvfuU5RFvc20A2ebLP3v4lo/5POa6vYc/kQ06YQ
GHx/pOpRfOae+2rz7x7n4VXXYmKf4VfdZV9EPV8SmFL5XoT33cPmOPSZY1kEyaumMqSWIgxm6a4s
v1Ow6YtH2ZdvNiDVDK0GUl315uUxqm9fJlmqZUZu1GaEbk+d3OwL0ItZ+OXK0LxufnMIPDUg8IV3
9kMEFrqvTFi/KWFEV85dWbjpNNEt5wUbNXt8FZ8q/qUTRSoypJW0bblNYM9tSBsD6FaEc15eZ/Tz
oq0SzXsT9LFHCrdlgy49AOArCZNhPxIVN4l44akxY95LvRAjb3giR03xw5HZDbUdr5S2PPoNMYm7
YDLi6Iihag2jz6HATvHAwko08h5DtPkQICG2oL8Du9g3TI/IB1xn9z4r+LBigeK74CtiVNbGD6fk
PftoC9ndua1OrnMndhBkOd7bQ9vySDuhsEZ8CTmwauProf5PZlLWr81x43zL9zP84CFnEZKJUhth
Gjfhp5/U1CG49Jlok4khTjJRJ1jtWfVSue/UuaMhCF5NLel1GAFw2ecwLiOmB98Uu+6LT+b1R81U
g8JxPXr98FloRXVTZgwBdh+ZNpSJLRoLjhcdYjTJY83oY6wL05tX8T9kLuTrtJyIgRJPoJ86itjM
CrwlQfVz/KRHVyYrl/t8g2o7XfiBkRrJEMJ54wl9eURsNXYvf4+Ievj01onz/DJMnyKkAvPIVs/P
D+7mKdXdIPcS62tyWzmdvhK9aGKX9NfP9Amdxjr50TAYCJxszuFtvD22MhSc4wrcfmZ8eprefvSb
GxVFUg4XJ/UxWja+T/o+Tl/V50ZJNQi92MBDKK01qGK5EiZfHuaobUmmWC0US6ZtgcE8MQ9lsuYv
hviqlw8MaZd+Zx+RcntmcJHWAHXF0IKa8t769mlT3P56cv4Rl30Mb6sLHAleAXTlZIXWvcsmMER0
HEyD3rvVUGxwurKnogIpclqKFQpAn6+P3EpBQUkkXw2HoRZCFjTl4DJoyX/W+ywVLWm1ESwhqICu
OwxfWcboUQRQBTEinl7VUbhAkEt2YTF1QFqboBG1RzZ88YDT5maLvlaN6PBkT6fzL6SvuXNBt/H/
Aab4qplCMxJSxeCi4QGnT7WKU1O/QwUxlAa4HRGqsAO2UsMB0IBAMcwPUCGsUz1t4kQOUV9S5GnN
5LH2ulpDJdHYoNgvMPiu8juOFN/Dyc2ii/NRV2nCv6jjz1ogKCKFo1yd7cwo1LydiY5BsS7MrQT5
ecAKTg6NA5Fpg4q+JNe/v7eBPPswYFUlvuKSSr1pqkDe0y1HUI9HzZF/WxEkdYEWC/6IRu6yZkuJ
4b1YViUaHh4ZJg6R/SVsTK4NYRBtJRAza+cftqPRbiXaLmdeHKlrdHsusZqrL60reG/UOE+Prp13
oKaddlOEzR6qcENZ+7TmBa1XVH9YvH+masqtT1mBky2X7fr7Mf6OZIsaHS7SUYKIdab/x0eGnBbO
h8Upe+xbVakkuj6DUIkj0/jqGrhtixNfpupKbZaAhy3yzxG7cYGfQVC96HdBP1eWbcZw/Ixh8sMl
Bu6Qj/gC41jAF0Fqcnjm+h9vHRMtrb7W/DucTQQKl6If6Tv1orFk5Vh7pY3dx3xgL7QGsqJX4xPz
GV7jSuC5qnbTkDyOBZvT/ASwgkyO4E7+4JCcZL/HvFis/51PHPBNVLV2USKv0xI7jz/87zb+IXIM
d7ZcLgsW6R/vl/z4AtAe7725owX6tnxlZt53KP9n9WLgzEuO50EAHSdda/fQPLPl5WrHdqKLB+QI
3OC83qu1VU2pjIBr4W2j+qeUB94wUeGo4ZMdv2jyQfNGrp0p4YBG/HMfTSpMZeKj32lfqCyhs+5a
UkrpYw4Gxj3MCEyKWcmi/2Kamz1TmqNaj1/3YfhCKSaOv2ZRSGJl+aXWB6hZvRC6s+i7iazc9xLS
5m3mwff/9Q8sJEmTn/A5GyMYLD3SFIDG+dBWM1QziPk7w9mQ8IxDcKn0sqLNDzLy9OX0P7ehlFlT
IkKgBcuobC1H8aA/gO3194ntpmwHRqBhUiAWFYRkMoNAcQbRQ90+8EH1QNwDVztLnMCVX3lxJL/L
XdfxnnpsPN7pzCi3fUQDXcsL6FYbfCd2WQEAjNjMRLC10o4Z3sk3YZji3W8Y0lOm5mRneyK11p9k
yINjgCUmYAYUzvqMmE0DRw5baI5r+/mlRJRiEBt3pUAkg3LJZBiT3A6SWEFZ0yOmyGWA6dHZUzBg
qQg2MaE5v6TiOepKCDG2QJI9U9gJ/YpLJHqqIK/ScjGkSzlF/Ta5aPyZo5eAKFOtn5cEMabefr4h
wckulIHNfdt96qUUwRFyDHPWz+HvEowsnnfLQrDZuE2wHSWd4pM8lGulasn5CFVadk8gfF66bKDI
zb/ZdQTiZD9akI7t5PHtg3Gn8MCLvForOBQLJSrSQgvuCoYXKWcRJq9i9Wt3WFfSI+JsCZwdoVD8
SR8ziImnKBuo1h6M/t6e69JuW79ZiEKb/oAjWBmTlTMENNcyCCYKAlDwnIHLgXZhUbQXMORokjeK
KFRsMp8D6WvQ6az+78E7LUrHzNImUZqhhzcUk8EX9Nqi8oaDujxyBRBNIHwt0MUTQ3PFigDiaTqh
/HH1WI5QmFXlG+yx01v8OXb/HIAaiqX3CLQ8qjBFNLZOkyFakAznj0IMg9/QmU6scUbuUnEdTQpT
SVPNIRulDXMfuDZCNVc3kOKfBKcGDaBAOphjpHnMV9sg/AnNaxJmaxwqvl1jhzIJTKVrxgC54Wda
zd3UUTsHhviZ6n9+b5LClfGK7VunjoKKupQl0PAG3JyHAnhbbQ0+3NZxYUNhv1YqkwAomUbDYrOl
n97YRbCZBzszS+b+c1JdQoHTY14TVE8IyGgKFwwgLoR/oTdbZ62ylS/pbPQ4O7Ve75AeMUSPXuAQ
xwf1WADBsiq3i5dnX3gNVpPYlK3i+XkVTCH0CP+qDxdKLoJUXsIe6x6fy7pfH+uf1D/7dLJhhr7D
KuO6+tjI1hFx6SBthtAmsIgb0Mml50QyZLU0YQcnbD0lJW6wvRi2y0qL16Dwq95/5HDqZjzn3g5f
9cDX1QZZGT/lkOjyrLLOFv7k/cFjiPcWFXhCTa9kfGmOMMVKCPlRKCbDHxnIYxyi/TIZs9lNAXId
Gu/yvqwBwAcXAcTh5REmmd+POdgmthHGVDTbf64GKp7JzTSbMdz0rxk/bq9uNXOel8ukXTFXEUgD
rn8F31iICy9gqMGWhQSBAJVeNy/+vBL9qSooDrMAaj9nWDABM4ryOXXflY+2fbAGQqJE65g+PcDb
0cwFXVu9MqovLNTqakfc4iGys7g9S0U6zGsRsPUBOabih0q/2/glstenxkriB8KkmkGOaC9SRyNa
ykbYwXGKkuHHS2HqgBEnoGyEzzuJcgfZB4BnEj6HqUEGLP+skj6BukCML3idFQwaiE2p9o3Bi17f
YCcKRYC8mSNr83bd5MGy0KEf5UQE4qVr2MK/rhKaB7U6fMxnetRCwwznrUjf2KPiaRk6IZPv/gYl
SzVa4lx1Ja8uZ7v8G/jZhdtU3ztX2FsbBxsZ5Z0AagjrgLirLvkLR2Z3sA/WeJCI/7I9DwepuaOc
kkilfvRjEO7jD6LKSARU3W1CL6b6umY09qNyWZuB6z4o/l5Trv8105ixOkML2q8j+LgHVQTBWM3y
bs6QU/pBqZnCjJRgDLwNc3qYdp5hSOidqtxZ7T2FqeDD6Ipp894mYCxGJjwcoOVMeXDimuphh6qK
pV9IZFSqmlnyYUaB910rEJoFQt5zbyTj5RxsdcWyqIfeSvDiL2cEDmK7gwzJ54HZHf3oRYaPlpuW
oZXUeWtOIjDHPRx7H6eDqGWjHbkKLkpt0rPq3F7/0r8XTx+3GGschVCgHSO3aRKVz55ahNlfhvN2
xhXflkFn/1VTY4FVuVf99wAxfd7fgCLa2yxsCDaDoC9CRmprpoFtno48S/aZDOZHV/YAdGU2uPLf
V3u/bFvF63e/A3edf6J4iI4Dg4suwaYDNfYdEZLJZPh5oHi1tyXQWQhWoSTXzyF5mYJjh0S/n3x7
k7JfBQHcFtEP5mML082ZzP4KRgDn0vecu5ZsIWhLr+mZdXEiWwceSJxu8bqJpmpjQeZ/WCxwZTmK
bipRnNRO97/p8R14+3YlnIFO65TXc3pS8F2ZUNtxX/qRaAqpFe2OuMT7/dwUaY4XlQrf8hZQpErh
r/oofMlqwz0dGKhZliJRM5nr0PWFp3rqDSnVGRrFIyXIUv6Xj4wbi4JPJOZ1IBY5ZTYd5Vimu5z9
C/kJeuwXUGdX2LI3i+lZURACBoPDYdnhl2D0ln4FUp4gyqLqPC6iKSLJ6qfq2ofjjmCJz66bgvnx
QwEtKHJWpykGQPVtVU5NoSQdCJJ3TzcOJOOqZ2nZ1JiHxkjVo9M3Fvr4KDUqAsPxZ3AlhzYF3m/N
PFjjaKsBqfZq6C5lRu2Dg4fX2gqVDgyDCe+BUre3rHqpSigYlp2zf4PdPYjUt0VSKVyTvt5IBKbu
X5pQTybCrZ6kVd98Nbh+IYJTTmEOQIRPKTjA5yhdvN3m4t5JV3zCUzjhu3ZCWQm3dW3R3IZ1tkuz
JQUUy7bvKCGq2JP4aZXGwd4gjVbZPAP9bwgymRpexMc+7xZYwEe4WEp2TXbqsrVn6mobcLuxwMN4
1+AJzkQwh5yJ5WbsPULEwjfA4BHDW72S/9o+DTGBDjEFvlN85LYZt7AQkG3AQNzVKl9BhHmLRCrc
aQa9TIiBubWDSYSYgX1AlC0a4Zvbz9zlLcuG3x/loYSW6w3M3+DvTpjyTififvtnPh9GVhtd67tL
IMxKMuUKqOqvrDNLqHTP7XB7NZsJ+enbBI7Al/MRKA6RfyAtTT2m0mAwvfFjAXO8czoKe5BKU5uA
4WPTywDUkCpRjgOsjdGELn16sfBT+62ufkwTVOYjPqDOEVO4tmTi5UM6xEXRGYoRCAr1EY2OnVQO
QwUi3eOEnVYM50xW88wpT6ueNePRg9KlXLbZNOBqdlIbZzoyWrfzlAZVJ9lWSjenlU5oCKNJhqzJ
aDN3
`protect end_protected
