-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ISjxVsXj0l031erQV6wADeGBCEFjDvzYssw+9dwnC71Fx8SYsynFvzy93FyDVYPBypmbGjOK643U
BPDvegJ6W/eSdPjYv5PxW4q99lpQu4KtT+C+udy5LVbcxvqry9buX+26YagcVzTyiE7kUMv6GB2W
LotDhwBYET7O7MjpA6RDEK7y5dG+h5+6sOAg8yfi7T9XSGieRWHNu2yRHsMz0LQNehdPNA2kJINe
l+OfC/ZF8K++otDL9qlamHKfFg7MRx0JqnSTeYO0chZiPGt5rSIpa+4N+jIsDiQpeXpcssOtR2Fp
P41znzFFXPIn82PIYi3EMoGMrbp/bFupiDwb6g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5744)
`protect data_block
WAWO4wn2aFHhW6z0IEGbJyb4g8rJEitH/t6QQzG/siqQW9VEnrCV8Wil4gNzG1DgtsDfeJRbnWRp
FwO2cC0gxw2W8uwyqrvby5CuJ/LTmPS6+mB9tI3iUBlLvgQH2hm+FexhkZ3pKAn4vRATkQv+O7i+
pInknJpum3N07zzXdUn/gAd7P6RQqM/F/j9Admn1nS1EU5217AR/68xeD4mVJttijOXj9x3wNaYw
UjUvsMpBoOYsWGInHf++q+8nSbjDnjZoArFuVGDDBpEDpnLvgnDoCEEYDAWpJMFnT9JmwQFFbYI3
pOacOB5rWQCkM3vxulII/zUC0krmEuYycMWZzZhcmfSIYbtO7S4o2CmPON3SSEoe0CEimawpNM/O
ggvui/lSy1iwF93LRaQ/JJle90ePeqs0pUi3J7YORGPI4bjdK5bBkUF9y5/zuMn4RWyRI/XKhofx
q6AjM8xdbW8yDG5ZF92XufmYJtsK0+R/Glvhx1wLu3X8AwyXyVhXBfN+PQgfGIkmoGCZcCZnYs+N
fkNJsD2GX47y1TaBcSRgLxTg/hQdkUl8aIucomeHBK8iSxeeKy7XBhKOKncktwynk82WAso+AaDw
R2DQpUXlZFxoNWVUFxNL9blz/Ov//BTWNjvHcpCFKzUIldBJOKABNZpLhDD2RndsSirCQItsAIrl
LvLk/JAg3QQG9e7coqfku+/ptxXQ8r4vPCSY5ScpQI4t1RleJkhTVLxeOpBwk4nzCmeYxztyC+I6
yZ+BfOjGxp1a4Pu+2pVQ0vP0YxkfRNd8CJIA3lAYPVeb72pAL04QhyJpRIHzHY8ZThLMBrHH+5CM
wH4x0b+wt9TvRDgy2j1iVqqZa8nBJsvYvCPJNMY3nldGfQX+pAnwNCkDVCb6iFA/iTjLE0rRQ+cG
CXlOWqSfxvZGWxclDG+Gy6oa+4olqDW+vs67f/RglaslUbnxtcY6LKxFOXo0ZEhnFnFw9vg4ar2E
F7x/mwAFb/5EMS8uaxjDDRgCnSat+fXafa3zuaz5TC1+7Ozxfo13HjpWePNXq+dxTn4KE+AmUZ4+
fkgUhCDbWZsKHUQgeVzKrH+mcWGSjZEFhSwAyL4oLvxgRtBuKZmzYbzPA3yGM5BOluxCQWr+g1v7
fj9aYKCu9xszMVf5C+a9DfTEZJ9HP4KZf0x0aNc56dFy3wU2UNL0D8Od/iMPoVMvnACy5y6nal90
KjS5Q4uhZrJc92q2yvh7zFcGC80pNiNOmoDU6C4sEmZYtIHE0y/h+vx7L4UPNFGFfwMJWTod02H+
cd3yzoIenQfh5ucvBqN//Q6Uik/8Pkfdsje5/6JIT19y3Al2566LPVhR9pP28TFv+QCfv+NR/Rel
CLxLFVlntvnk3stJv3dlkKhQZsAqEwzJ1arwbMC+xYg4tTToO/NWSrC1Hj2jEvecSVYwtC+1KTDt
RGiWl6+x7OMvZcrEa6AgoPi/y+n7X+VKUaPGTQfDmavesheuuNZ1xNOTG+xT7LRh0obDnAyWkZ0a
awOj4g+Ar3no/fP58q1JyhUZ90m/nbh2Ah1R6jlgD68lWdu8mkLZ8PTEWCfQfLifW9QaVIp6a3HC
25ia0pg7HgNvq+6hIYStPEl+9kQc2AGPQBbGmMswgJCtr1XRn83zR1T9xBBL4nTXXZ7IIL9JSWhP
KD3azMTu7sAjqOKs4hVe3O8lXkLZRW6Lo1daFzXIe1JaX0ESm35r75nlwcY2ec9wY6nUX4e7ZDhM
daibD0FIhtSk4yvOWt/a+SnpIbT6dlspUbUnBKq0MmKIK9m0gQa8MtqJLLcXJ8jFvPuJKhQh90tG
UQD8+VOFzbsRu0YSWKx5dm/tAbqQXaxqGt5Cr6oRIB5tOmYxBV3TibUWROOrMaVMbH3QsYYQNnWB
wRKTec/v7I/SNg/qfmpgjrOzHLbL48OXy5VjWrXbmcRW04GS/HSbhKNZUfIwW3+ki+4O1fGkmwd2
nqNpcxtPLwevzWCKYH7TK+83IOszqEpuHeuvC4NRANsnXYZsjKiFxt/5MkcOvRk7B2mfFf2klNsa
TnM8DsVaIpVjU2p1nxOy0WIjK6mh2ExHUNcyuHwuLsQcT0L7GdAWZharvof+JNkenu9iYmx756Sd
/+tG3h4SptJBfVp5wVsrqbm6XakzFz4nhsocpi1jNPKLMwzIpqN5K6m4xFL7l4z958dMBmjbIxMv
p6KcOQsHFeqyYwNWglxoo30Nmaq0pt2PoqflNE+eTRkQ/FzqpjYyepAp5kmS/e8uTKERlMEa0TbO
3Is0XmkA8aLlf8TgafLSxjAFd+MpHTrD2twE2LFK6+cfYm1X55/zauVYaEahuDhSy/NrvM1nEac8
xI0UEJV4PB73iyPpWYJj+EaaSfewkx2kU5NAnieO62ujSjHnt2DkyKJlQhkV5lN26+DmZcRDO7bx
/KZPJKzcKW1+LNsZ9ac6WpGoqnkpDsGA9XECR2HS5oCPPra1b0UHJuSbP37zO0wL24raXWksDDSF
CAHPPC/HvvH6wt5aMieh36IxuB/ru5LrWMd+wiGIHoqB9sRocXnob5tpqb9c/m7bNPdenf6rAPUv
vwC7QVZfRDw+0LZmFZk21RkNQKOrc6b3HyPTCRFjRvN94pKjIlFpBzIp+V2S8SQva4GmG8aGi+hy
LfINKusnme0cgLsNi97J1yDAc3y3AknSw9OXmTKpf2oyNC62PT1V3/TRzxVyu5XpcxQNt49we085
4ybnG0JMeYVhbD2MF5rukMBjAYxJXI1Hpf5X5igt5SBg23uXq2GN83iUPVLRK1V741tjNAKij0V8
43rLEYfp1EM/OGx8kddW3Em+dyS8gD6k21xxKZtNrOglRhtBrv76zhZky48/y7sgSomzeiu/eiYr
NyrDts616V34YD9M1tqNvmC98kfjg429dZBxgtdwfzxNWDMW4e3oy7k/PEAvwN04j3vMjJa+011z
ZECbcZQxKRWh26pflwf2v3fkfYHlmfqXC6jXAAy8o66aZGsj909TTtklP8hI4O83tpqByF7FIetI
DZYs4pE7FBPM6h7QolNbzFnauQlrMLGE5eNAddHfTgApkzlw7R/b7js6dHLEM0qYBN5nptBzQrM5
OlFIL97npw76XNrGEBiT+1H1iuO4o/PAQ35FQtSHFmGhh6wXqKldIP1FaEXtbhgEHq6n0c5zyMm6
KStyVCLInhJDlrrEqmWGpORVaGN9rf8etxW4yIFpDsAKnmqBkP/If1o820sfwmQwWi3E0MzGLC81
N5HeE89P0tMO9LhBYKHyzZ6ZuhrCJNI3RcUd3n6UIsy2c9WiStquEt/CA5CX18Ys0/X8F1zh9RCB
+TLBaSe+VZ1EHJYLpaOLAH+9FPjeqdb8PiRMsuU/iAmjuJKsMDxeQffSTGHpwa7p2VVUgXTpFb1e
l1icloS7T09BkL+qAN8a04N5472C6uA3f2gGUbM6MBJ8yCyMvkU8XO3/V2wR6Kw+MBOvAP8IdxQ8
rYUbFmZshMRxTmTAarVeailHqRHxpe1BqVcdL1K/iFp4weuMIVECHLply7cz5dOSxGhXf082FlQW
I4cZpOsRER45P3/fPKQ/lwpJM4moxXYTBPFGGipE21hvju/VPH0zb4tsiyCLpi8+JtSMjUPW78Qy
UZkXkHprLL062fUlZLy91Guhckixu3RQ4Mu4PcqpeHpC7YyezBfMalg+qEVtkdbZeEKp8GRG/H6i
btyp0yNHojx6LNHdDrh0kCEC0nK9E/UcrSc44bRXpGZWzii7CThaJW89R124ZHTf8bqrj1iSvbrV
0hx7Mc47TqGuBY+Dl/tr3JdPwMTMQLUHEWiBeYzudif4E/vU2s6Y3oFJwKhv6kXSsJYPdzfvvse3
5oUgtnnsEwEcjrBH4reU/cJH7S9CNFLTdM5IBY+t+3bJaZB5sgpLfJq7iUYRJOjVee7zq34X6Dgh
A+BUKHQczSHEHD8payXBaLXGO/a+vu9NJcL9hhixbZEgICXkuGDJMln0VqyXWHVomjoCYYSRgdgg
bk6DmkW6kFhXH21gUtrUNStXCPOCf6tnox/6Werk7CPjENMnIpWOEIJj8g6+JVdGu5VkWSlCoiXn
J8x51gxSitcJ9vmdU8AYpCXa/XJ7t6wUIk8E1NaCLFZU4XrLni9aOj0qNHi+a4cQle5emS9VoqSl
Hm7vR1rQHH2hIyP4c8m16GhOS05AuOjz19+pDbj7ORdmREjQMNZ3LPY4QsMpG1Jmkc5rlIEIL+24
0onNQwBZ0NoV6tSCZn7xNETY0plEf4tv4JfHib50KE+BNQ/TozcpMVcfOClKo9Dk5PTmk3HVMeMq
gGZcuNcvp5lR1uun/pdmEZ9qjSSdRDLh+tZvsY7jtz1IGABm4M6pXFExk6K3JSpUMq8ILvAYIjjj
H2YiaQtrnj2OCNJws0JlkoEok11u3OMLF82YX3Qfu0yFti+gQUaiLJlR8hUZnpRALv8sv4Ywunmv
RkcnFzXfSy+/z70hvWF80IhNYPGG62jpScxP1YRamgsiHiK4PCK9tMsBSmhNUjdkZk5bXK0iLoI/
tNvosiYShPVrjqXziSAryk+cEI5Ghf28FMTP/uoadhWbOdCjvJdAbqSjRGsh5UKbunpMZJn6ftnI
DAf+UOxS8gW6lxFvWdGTWxOKekHNufARHo4Uv3+WXLjuHlTPdaDa4ZXQV4bYvnpbQb8tRTLx5SEj
sekhzGx7XgLJrChuOgEtQiIuyAC9Gvz9MSjB/hqgomOpUUPAlnocjkZ//R1bZ+p+5ZsbwzkZvw0F
GlentNIk4mLWjw2VqjoLVtWe5ebrt3qahmKuth5cAkCHGYEBb84TYLF5epqsVNr7dd8oPMPTAcnt
i1BiyTXrdGjtPllI7wefShoypVYDodNWkkY+qXl6ywwfCen7A6Q+tu5bpBOW9lvxQnQsowLdZd5C
DcJePCS0vi8U8jASsMJuziWNIksWu0lrF3042vufIvCRvnHW8NDUIMLBLALUd7rqNmhgxB9/jh4a
y7AiQdJNVEzMfSz1sIydwvPyCKy1zF5DqUlnWxzEr4S0flDz53t/fpNcPHBmJpb67DKZCoDBQKD+
V20l7faG27+YJ9bGCc+MZIlg7JWQib96m7BzncE1J+Oi9XtgmNaFJfXzsRjpaQF8aGcXIR8l1Uvr
rr1Yqt0BdE7lonuJnQR1YYg5LAyVCTanISOBN1SY293vNONPd16SOwtf/b+2oAeLfdC6/KbHS3as
ygLNZPb8TIq5T/EYwCkjvR4xACMAKB/QbGMQNEWknTy8u93kdsRrePf4FwaJUG0c2i11jolAqPi5
bZQNhh9yzLHAUKk/S/PrxkL//NH0qngjTG79VEOhE+MivPTpKJKv36Wk37WoIOUJ71Y1LlVtEed9
A56PwWi1aVs+zh7Gj/DB41hh//bh5Ehem9LTGFqUwyg6HwQa/rxhLycIQhhzKK/w2Qul/Ex9pVoC
D6dgjc771hULKBlwEnRkgKUCUsk182KIyk+g14ZIQe4wAR9zCICop5viQc6QgUcisXJJtRkP8t9m
5MMVpD/lPPPIcfkKcb1mbmwdDu/u0uyzMxIun2U+5Y43uD1i53MiUTg0v2g3ItMoewNtzr0M4Ybj
b1pkRdPYf3lASiGF+IWLIJX+fyPlH1DzsJy+AXj575e4gFKEubX+H5XtSkLwjN7bWo0K+PtnAo66
q1selmLAjt+kQ7nDzEmWgo74ht+mCJuyvikBuzQBMkG44HUF6yaIWqG5h+j5WIPnw2mR7PXVXCzV
g53OXUz+lDg8jc0romtdYnE8R9Hp+8wTHewqGjINIcuTdNbZWD0jl51rhNf32fgAy6NQ6uE8Tru4
IgLDmMSwQhRcJUdjqMiAJ/SRZCLoZgBdj5pajI1nc0NTpcgkJzrZbZdwFjJdiS14+nAF4byXt4sU
xFloo9mCDsF4ohMcHhj9zeWEGnON7M1fhhRkPo4GufBSYN096Wn3HokJJVWVU2FVY5TPaH3ACVN5
96Kk+kJd3S9dZ5uQnGxjZ26WXWGGmM/VwtCv3u6J1hSbXSHUsl8Q7vPsqiVJlW6oPEU0Y5U7KmO5
C0ZrKbWjBKHR+n9KGl4NSH7oAuICuxTdZ54XlWHYj2OryfG+IPb8x0lwHOeqwGe+WdAbG7DhEvFJ
ctwpZVFow4ep19/ghL+ZzEXkHsDgPdMinylN9uIr7rLjgXUIH/c+QQJ+uyDtC3azLfKeg621Fgsp
5JeN8QntkY1Yu1V4bKagiNWcAwzwLRuGQPCCWohXxGMEblhXLIYPvtB68fyiu6Dkw4OmUCheNBOB
a+0AQufJmB2uNJUBcN+9+O8220ZS2cwCjML1LS3w2VdZristNaIv+J30OxPx9BhfZvs5Tc5cymM5
EwZ428d4rbm2E6D7yL+L3U9MGmEUY+GV8EuRjxYxxrFx+zA0k4pfEPk2sps8C+Fw1iqQ6DPkEkz7
BRzkx+NjqpJpjHEW50uOqEuM5U2xPKe0mCEjAkJ5R0gCLwWzANFTmeNa8NxMqXmBxjjXL7CUX5bf
m25tlXafphG9d88TeUdoREKmEP8EC5+ZngS3yZZ9zTZ5A4sykzO0eax73mgGMqxEnn5owY5lD3Pz
IkiQWdOb+bj74Cq2ZR3/J/MLEiNnd8bLOI1aGLP6RIdwCnUSKQf7UwaxB9j6pYwlcnCFFJh67WTB
EFaDymyFGZx38Rs52GSkCfRe8W48jVVe9OHprXsCRBCUXd4OEgJ8TT3piQqCMDhS99RnIPodF+yG
VPsgc3dHA0Tchxc74xKvgMGA3KZm1uAY7mTln9xGLm0hKlYahvZFX6Qo9DKtR4mFBHSrsVPmfknQ
xDD3iEoj5CgACS/lAfSoRyFvUtLY6Fu7bubSHyRtY9IhMvgDk7xwXSMpkpgbVitJRd2D7TFBtbXO
XZ1XUSC58bYFHbq78g2DYiW0QIxRImwLzQ2UQQK49VcBYwDjH8dK2Rh1/4I4aH56emmHfvqjWuou
AH0arJgfSEe+m0Iu+OMVid5k6DdYdCZpABtkJnpk57OqPiN50uGTXtcqRLaDmawZoDn4WOSTepAL
TWgaRs058VXui+0S8rfB7teHAQR9r+zd6WMCIV0D4y2Aw9DITx5jPEdI7VBAohsQCMgJRqWO2NWs
60wmnpvrUEROueDCENapbaVDUWq43A1vFAew1DRtj/kvsGhEW7JcHQ1umYIcV+tuMDHMzeqV372d
pavzaTx44rSG3q7VWjw76lnARLUC6FOMO+a3MrCRXNvbJyUeWy6I8M2CMe+PTaamLXZEhHiwVSUZ
GwzWnezu5TtUxoZnjbGaBSc3hK7iuMUPIB2501mTfdmbhC74Cb/iIq+e8je7DoEUOauharadBKcs
WU6XzvgkLFGYIP9dPg4mc4K597X2bYFJcVvg9BM6XRwZSEi8aEh+mBkhuZwY/o7Rq/xG6qBWZK3P
E48C9ws2ioJfcdOMmAMLZ/Cbgqf69rE3JOfajfrBSKOCc5Yy1pPn1Or/gQ2MMCg8fNCGWsjkcE2c
OXPWx7pbLr+8VOsJ4ZnCvcb3doxT4juyLLPmxlQJjGsbgklHlLE7xNll/yKbkF2gXv15KUkx/D6T
ulX7fnXwvw3528G8UIRQ0/Ad58YYSzeA+CeN8bjUouxR2+7dUWeyFHICLbU=
`protect end_protected
