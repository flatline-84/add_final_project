-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
V8bvM7/fY5fiL8NPtxZSLsbF2HctXISZtBapGfEjiONzXNAhBJIHTHpWB/1ft9Yjt5pVHkZJYdNV
rrx6VGaIVS5S4eMJSfu74UaQQr3ypeEIj2tlP57WW0ccgGEeWW72cHD+gj4qUwIQNIOzvajcLSba
qNX+gEqALz68Pkv6Cw9VHSevke1r3iQzQmObZyMg5+pNBSFwKbZTpmmXUsciBNQEV+22PDD5Tsqs
/2nuyX+6t7nATl+ZQxgjVAL+hqIa0yn1xF/QFmT3KmHOiuLpoewReBm4vv7go2tpZ/EY7EScMqL7
nQcUZq5HhjGsroI6ILjJeEw3ltNOfUrN1IFDxw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10336)
`protect data_block
ObiGYRYFpUkwB647/MVZUTGsNSOCG24cFdJxJ0MSUpdE2hOzLWsfkCOEfKWyEcUHv33MLTuB7fxd
lkozn+D5x7ucGceqGxKdkpsq856yoJi2yiZKt9vrjsybHPwgDQkpG6oFsRLvIxXueOSPA17lKECU
1WYLwd/3VXq3oms05YisxQ1Fo7/n2TRMXoqI9sJjMvZwv92KAfSrQ9CLtpJg8kALT/ud+BNgatbs
dsduJe5Kggy7EVEDQzZwfv1PDjjPKMeQ6/b5+jS9j8WbeT8/EDb02CAr7h0VXb91teuclbl4Q2q8
VtXsAl/M8BMxQKe+B6ThQT/GKOLFKleh3peQ/SJwylZfi0BVvqCBoyH9yWxlqD4jPwFemv5N2jtw
geGBYoL+5h7mXt6q9ZJz+utF7B8hh/WsvqWf76M4nHLaGJUZxYsYGxb0zMUutcZWI/mqfJ8kZnx8
dVp2k4Fm0D/x0U0d10Qt1C6PfKPAvGmtDBj7p3QTWFsYhuEGLFmRYpwveGrA3nBtGy7pEMQmp0A9
yh8vaoS4JbnYgnM2KOxXHNycBVtKJULL6LRXVe3WG1vbwAcZ8iKlbzSCzwMiI8RN7NMAQvvv6kwQ
+/ud0UxrpDirtxNYCr6ON8ygokhGDs5xGmWCUX7/+YN7A4+Naxc3VdqjD5REKdJzjcA2ezVI3F0o
5i/sm9x0J7nDLNKzxRaccw92daG9BB6e3NULI9yz6VOkeJBu8yrIQphT/l6PQMzmjZXI7o+01fI6
EUKVBX68vCBIgq96OIZsGe1SaTH3vaS7OKFY2SYFt/6IKTP1f/hBFp5ORAIkkOcxo9i6lEvcCf1A
w6AZwk6kXXtPO8GTbYGTsA7IPhQtzBJQHl7h1C+5QPRNMmtPlGsmnx3lMoNggipcCKQMiXcdjdQ+
SF8uNo5xpAr+9SOYdCgWOg3kknDboXmRMT0U33ixuWg723txzguEet8LxyGdA/ue/eUazhFF6ihn
cyjf99DDb8ceO6BCLLgfo2Ql6cNSdcDJ1bFx5DDlVYT1dvgmp7QrQEm2RWv1s3lYSmqILeqF2Xez
S78LRo5KEheooJa4apCQHITB0nC+Y/Lep6g17n7yINJIf/gMzdYhhSMcunmuU1iZCSAsvxnBli2F
t3SPJGtg3a+cGEJyubzkELSuelLd7OkxuyesNWmw+AFO6s3kHNPr91Dl2zcTmHhCHMIQvh+al+iE
BByW8ShkiHMPOLDFCUDwq5JJ4V/9ph6Z0rfjZHN/MZ3AUtBBUES4s/Oa6DqD8ZN0m4NynjUxkDOl
aNf6AUifK9xcdq1poQ2zyJ/TTd9HvKufROJc/3Hz9uS1ROlKLFDY37M/4wKk7r4Cli5zfoiqBtpG
y9LqEwsqiOVeS5V/UzWKHy0pb3YPgmUyCrFnJLOKb05Yu5PjhXZDjbE4Wbn8d0dAIFFkyAFVXHSL
SOWsNTYq5OyKn1xLBNydhpXb60zc77XlbGGXWg4E4e+AvJU9WcBxQIOe4/aY4JC8YzbXUU/Hfcvr
N8JSXjj/EJEJ1t8PwVKIgfCY3CblhJjWSaOPlCHziXn0W47UPEGTrRhL3k2OUNlyFA2F3odB000J
8cFaYlTJN0ullibuvp8gRewXrohQd8ehnYkH0oC/DgUQzV5VyAbIjTKDJeM3STz6GuZCXAGuGPFU
lakmy3nOj0q5uitgJcdPOTmTZ4oxyDNkWhKuTBiyMD0u6PMDgN/l3AodZ4mw8iMdvhbLMN7kPH/7
Tqfoa1ZDFoSjwZDRllu3LtWD6KfzvXm1MLu3w5wMMXrlWLniUy+lb7WTron2A7Td6E5VGdGUEFvs
QP7D373KgsVE0M05Y9+76rYMeGCDC+NJSBvSqNY/lfV2boXKt3C48WKM+6ihfrqwmr9j/abKKjyl
jPj1efs5KPGP0yEfpoDkk4XpgTRRqduWwfhUL0vHci+Ez4sVeAMhs3KApPw10g8FuFnyGSKTvuc3
ZyHpVnuUirbx6Nmfh0DOBfdGp+M4gkO5efsF7qsnZ6nspIYOqJfg0dLSJVMms0ODVApSaGZRhgKJ
bhHZ7s7ikJ/l8EU1De5B/Wi8Vq7rIQaMqur/tY6U9u1PoWbwmWwCIBQCuHAj5NJgubYebnoo2tIg
sOxueQvz9jhNWnoc0NDzf8PahTq529xDCBd2z13qLDh0+2Swd8kMZ1EIJzVOg2yKDpthKdKw4Ibw
q2zKI+akR8cwcxZzbAdHmIAMd8qG7aiYqsa9+gsmnPKOwY8dUFp93UF8CPHrs0z+/G2G5hXgxEoB
xY6c5lCBfBNQ0xgIwXiKKrWK3y6ksJ4hcopgVHVTr3nrq7f22Kqb5HWFIVRcWh9UPZFnaxRSoObO
3K4Cv1K3rnPBpnxkgPF3JBko7c4IY7K80gYimOQMADHSQnOpzfuE83Wxksbqspj33ul35LNY9rcF
D0EKhEFq89xlm3iuFGif5SkH4p76uVqEBIULfdXniMxtBXiJouBlyWRhEX1MoXH4LM/KExZREkTa
DiVfM1IKZdu500juVXjUApvEOgsNt0NjyuwOahzF4/uYOCQuVXnKG3IISIvJc393wNL8yb6ihfhE
jEjVwVVZzRNqULVW/3UEYU20i+71Z+XKOm7b8wFMV3ATAGY1JBm1jFRNNCTpAnegoHGEujRc09Qb
d6IGIkpfwpZpafCdMN3QvKtPLEHGmR3UgjWj0n6xl9jvFC9i6Y8gibljFEUM7wqZjQv6P1tlITez
nByhbgdtSbV+kUucPOCig8TJxHlRauFVJ9v41jo3Ag0lLLpPqbXckOayj4gX28ObjPubAN+R5hFD
2kJsVnsS5WF4mWOrYFoBTaZEBEbvzj3LFMFa4gSKuuC54aGVlqFEkUzzVO3aosu8E38CzBRIXkgv
7/2nK/c98rjfpFbpLvLuir9898GAQoKvxExNzU+5+0T+ki7XWQSGZdRRStOL56yMdqtGPPGxxupo
30S23iuirrFz6Q0FacwNmTgS9R/K4oJeRJlOejDVnxNYZvGqvxV8doFFhxiDkEUjzB4Rd6UDdpPI
u+eX852VIhs5tmhncQ8qIFDVZxmwww1VdzEjg47DOhlbUr/tB5vSDl+HaWWWqP1OOPZgu50MViuX
h1QqJq9CYUYaKFlBNAxAUb7c23q72M6UmwIfHC0YIbJrxo+osTpeMx9ca96BLnPu0LWbA80vO+Wa
4R6w5FUIJei7V6CyAAddf5ysrtoaCbV5jaAVocvriWiZQQ+5hShp4ITlyQr1CFZlSMaZ7t8Ok5q5
uVobh1GQq2pKrlajHZHnzbxxGV0Qx2rRoy7BOgsoPz+74YGWPxona6zrK02xfkPYpthCCoVNeyTZ
zN6QdlafFAHo710Hk83wr4jmwXLYLAe1DEYBAPAEGvYec/G0c3Ue2RuAxRBovdX718p2IQOJwFSj
Nt5XszsrjvDwBcvQjlJofOAaPgI2oDN+bef+Suza88Rz863ga/MqPgsJ19WVXggMJkv0F91hrjGk
S8px7EyMWdLJqRjLGTgjTcorfBdoxBNSG8Ir9lRgKQutkzxkJpzYlFuRTf4wEseJmwD7DYDdW/i3
YQxnJ3HciqoG4IpkzuPHDGIqlp790fSZbSgQjlHGPIuSUxqxVC/u197/kltuQcfY4PKQT9E9sIvq
fHG+zwywChsQ2x5vOgrEq/ye731G4M9XnckzUkYidw/RLtsoD60zhYJWwFDaEEtcyZcXc5aS9azp
oxTkY/7TgP1n6Jgh+V+NL/YqNkqWtp5hT8tDfTBZ/Zn+6egrwE2UdtLbmVTg0qsVcVDZNLA/arCI
NEeFgMl2bqmQLjsIS4xrjtE2iPQxlANvGPMrzjV9mGLca+9YfPi7XwWCXpCzxFL4w91QnduDI3mm
hg5wNBg1ISp0qbD3c++kIHOsb3sWN+ffPBDNpZLco5JaUbghPUaua5+2fWD2DALMfQhZ7GIyokbZ
AuGQwwfsM3tt+QMOe3C5GelNEi/Zgf7Cl9i+jRrNmGvG6lCLXkXfk+PCht+DkSUAdtfut5IGWLpP
JRLcxhSZbyVjeEK3UQ1plUDmjch4zSric3nKW7yjsxQdwYkSieONxRnkpwffHETfpxdXHFZm++f0
9AwCM6A5JEajM5wp9Y4BwY49hOxrFuH/yygqK3F9BZer+qaRWfLro4BjEkv/SqJ3nXut6w3ums2I
6xrpypExe0ZDY4HyL/3FWQJd0mPYClIrn9bSzpObGHg/GK0t68XVhgcC6F4sUads0R6F6NzKTs66
DSUMYQsC07nlD6Sf02NfMo0+egzpDM9HY4XKGFg8rFbQ1+PO937JVzGfnutFF4gVZ+/Y5t0G129c
iE4U56sM+RvqbpTQaSIIHj79cnQ0E6sPuTN+5oR8F1DGhRfa5cSw8IuFp2VROhwitQ7yEuRTQwVR
E2RuqvdqwvaRa0tTa1Yj4re5dGocNnSz45SHIaaN98V6YGJkyOO7yUq/K/GDOo2LJD/ZJNOznu3q
tV6qoAU1hBMK3806aCwzXWUlrRWCWYNLKdqLOw/VGNIR/vivrw+sI6W0ZnumAKHMtIvRiN/RXF0b
o64k8baKuemL4kUdtN7f+N1RQSpaO2Me40PwSsE1q9kl3LoH+C9xuCNxSUzy6gETq4z38iO1kBy2
ZwZ6nM4/jdY5zGhG3/D/9rDyL7kBpTCbBmvwbUO2iaxWbSPycruaomWXAB+dnbo0FpP9x0mNlvXK
Z6wjxeZw4h1dxVhpX9LshZlIY72AWN9nOwuWO1P531/T0n5e7gXC51eqjQkJoZsW59C8ormM1xT2
GCmmbPgezBGNJBUXl2HMAnMo6akhcmC8PXUkBpabzp5qjRmtaJEnme2ed/i5pXXtWMtEhJrXzl+i
PU+cDn7IBXuBV1/vpoZ7K7G/1exF3AoDioxb3A+j5sRSHq/Ya2jFkOcurywo/SvAx8e53s5WekSc
np+4lkj3Y6/GY/dt7ZfoDoLwzSNiYx+XGXbKmVarWZsyvk2GqQpqdeIf8AaI22PFHywJiN2YY2SD
UNR/eTZ1nNMxFl8gf04nuYZFRdPLOfpF6MkNaTwGb69Sm1fZraP0SqKxPegDsDMpwRXEFtCTJd3K
slO5TbOh0OtZ0bI65VBvKAXg3wCG8hENxCL+2IrlF5EHtU/1QXJMc6X1XnF3sabEwfezn2zzf7er
2JwbzQ4y1z3BWJGzVa4UwoEzoQ9IRltUDLgyiJU5eXwvCHQQ3bF1zV5euQfXRf+G3QjgbhPXA1Cv
ZIP6M7GFjYgeFXB/Wbtgq7Fot0Pm9E2j9lUVOW9VjKamZz0pavhAKO6qCfTxo53RNY8QLGYsrPeo
y7nHaUMt9oep0Z6W62AwYnbrMEXk2tjMq5fYoU2Yyfqo1jYktD23QxgZIF+bnEMJNw2/bbOGrdq/
9Ibd4bzODMdvYIUEXtodNUtonfUyddPuCUqTtPsizoRmndOCBHNUmYKw/7gCym66v3ywUsY48nFn
NiKwLDhI9daaEarSbKhO0HZFLG3vU8CyKQTop4Zejt0n6/6yMtOjerI5HJIUP8B4BpugYzU2oNPF
XtjW1x0W1Clrt6blxsldYC8Cf8Uvl+ZscluMGt2Vn3RE3DoouoobhoSEudZr79th9PcIz8SwT1+V
Dc3jv98yF6qTZzGbcdB9kVUq+B7SpoWxUOL3jQiM/UabfBXV1Mkku0ctDS87xublk/8UpYdivbRW
r3mAy2PzlNhefl0KuZkfEr/rEkCTpuX++lAlyC9ClzgTo5hzpLvvzGtLCgsZ9IbkvskZE8v6sR7D
EQQNvIQKOFMfYQqBRuVvzZ4egWlEoYxJOhzPAohRHPhohv4CGVBI2oBwBJn3VmZOE5SFFbjZSYQF
bh1IOhB2fDPQ9Jbx/zUycjShmjwLDD2N8JFFXMWF4T3gQkFPeVhaxv4twyGGDp2X5bQa/h0tjeyX
ivxBr+yPRRK8tMgmaxZLommxXna5FRHKNGseux0yGCn0d/S+YNIfMkTnzsT1+QDoo130hHJTa+nA
I5cMYTVAPlBqwYVfEPn1PL2iNCDrYBobSP16RG65TFBHCe4Jk8tq6snbuW7EANttMInBbmp7TvqY
S2SH5fmUTz7WNLcBbiZFrc/wye+4oNjlT098v/50KKBnuRadStEs+zNN9v7d7CF0oQnJEU5aS8Tv
h/pJmQpqVt8mitAF/T5MKBe9DMYNpHS5YmyfGjLHBMtvLw2mkw8Fep93nFkggvQ1c2ld9xlsWfkx
MDki+yeiCNNyH87vLZxqMpocSChNR3LbTcM5ERtUFVwxqd/dxgBw6J4aPchi/YLYGHD/XJUTCR0P
9xGIeJ4HBgWs3KZb+6IfBBYk1LCStyHZnMEg95ytG0fLzDigV2KF/BjWfInfp2TLCSa73d3SlwlA
XQvEi8FW/cvaIkEbQ3RprOQAKcvjsxq9y9ehjvanai9/PGzxpJTYSafNuQeQNYl1VZgc97iEttip
3/DhuGU9znAv30Ep96uDZVfS2Z7a3h2zjzPXiRS0SYDK8HVebJVPt0qVQXq/zgz05bGQUvPcLSqV
ZTFZWWUGulLYxxBqs6SCm+ngAIIdYhWJIfn+MkBDn4kEsZ/cmbBN5PtO9Y2qSx0Psv+gKf0Pl5gr
bJWhlxbLcx1bJC2uLcj7DGEqCaM3XpgzwrcpoysDULc4lcoN/w6Ub6I45Ntul9HdqXC3z7bSpF0h
Ck9TGa2pmWesO2/h8+2gmMBM8YS18bgPQ7TRKS/SbYdRvfk/jRZ5xgTYJU9me/YfeNbo6QkzXTk1
yT0rSKN7wJORX8lQgXTq5+ITCwda7fo95+OUbqpyGRkiVCksX41cWfSP8xmlOO2OVwUK4KxrOosX
K0z3yo4cL59FXU3KivFvVsfaPuY2fdaxUEA5ZKAhxS9QOlQo9mvwfwAoqJZOGkjsTX2RPWzCXK6+
gIpolJILthMc6bq4694BdX7Zd/gGC4fpnkzkrRT8Q7+osSNAquWZhecy87KNT1NcsJsJmvToVHnL
bL1vQgguGi9izNkruxRQ+/JHqQoltjQksPpLzHeh9PU3sUfqD8tAyb+cjTUzUDBi4T/0WsEM+JI0
XqxKAoPnT/M2Txsa6YX0rG5T4aWftcx1R5kG9T0mKRYhH1QmpZLNljJGZf3siHeGkL9g9V0lqVWW
fNL/fBYp5CF44xpbRm+Bd/Y8hIonNvA0Au9EpzQKJAinQyBtKkGFEMmMGLTfCOVMt7XVwtngvZda
mr99hPUmckTWeR6Wi/FvwIAWPXSawjWYrA6e8RHvv3VIBUO8sTSwk2uDi8uBbSxGHrI9Tjz833Ht
IcU9I1CTmp+Flbp4k6eSo4Wq+L/JV72hEwCCEb1LmB2m0BhSAhNf7kS+X1Y3vrisLzkdw1uE+NOE
IrNGuesq4aACzr0GzglL260+vdgPW0BYQU8Pa52XCUD8k9prGRtN4YtzJsBTl57ZWz2erPa/tn9r
a80CorvVbBpOtFot/uHqxfBGtW9d1CT7jnCnV6tLW8GJCG4s6c50HV5pwYVXhrxDm1M2l5oXpyM9
C8ZxfVVwYt4PQYuDFF8cpjB8fuZj2+ItKI5dAD+mWV/T38gJkI/b2YP6HsfHcNNFaitJWwZNYR8d
0s7meZqSV07Y1dyX3Fn/X2C1yOX3rOQMmSJLql4r6Y6O7+bHuJDqx2WlFbuGeMYRadZAycLhAplb
qWeLUhdgZTjXXt6lWgXjmWdNIHDU+bAVb0Ue4FBYIbtN+C5VCnuPqGiARskWXVMx3m6y5mUYWWgL
LbOnxAR5Kk5Qwk7eEXRot4R13WZweGVqJPnYlwa2erEGEhSMmk/rSR36gW/wQFwEhjHP28/fZ5CS
g1s8taK+hUFoKMpZttXqvB1OOZIOwz7+rb5HFWb6EVflGbYpl3qFZfyJpIJ5XA1oTzLwfMIDjGiF
VqpD+hXzsAp/owqDWd5xLSuo4V7pDFHb4/BVZMdu/IeqcWT98yqTPooD7T0cj7sPmWDsPuqdMn2C
Jop3vq/IuSgrPY00lxB5zBYugWr0+3qmW0Da+vVvQzcPUPgyGdyCOycO4Nc7yW5n3871rvHLJm9g
4NPLST17rFTIwyiN3MImH8rlI2eTddsMdKU0HwQLnQt+RjoHxxfmvvi1vOfaRWkk8cobLv3UDETN
btZrH1AHD4hk4Qsj4n7UY0cNYhQOnaMuKSEHE8+5kh9TTYgtZCx87DJwooSJetAu/uPOyBdflSAs
YRcwAbPd6/fLDgg/57M9LmuZ0LiPiLKs+1gSSLEul/HiH9Uu9k0NYpoDQN/IoN4dKMeOchVHGTrA
c23zi2yRg0x104R+YLQs5ZH9p7CADfgl1IIJ8O92xupLcoKI7TRNOcL+f5c/dIS86eZjPSMKSsRa
Sz7bDrOeefxrSnorEyKqQHb8Mv/nFD1ahve/4FnVqRkt0QvAuXtVtW+hqg90ED4f5qZp/GTSpTAo
19KdfYoD+L6845vUT70eJtKqDS0BRmGO+Zfm2y8BXaGQGs/BX+vlbSXPajaX3N6w/C89npMzCJf0
3KLAv6m/uGFeKN06+lF1T6YKFspzLO+UZdtrZ6WVuJpfx+zz3ULOnfg+5Zdg3ODs+iUXWgrtpIV1
gLO3eJ0UFl18fOVs+csH7srK7VCUvlCnyKJ+IXGXtaGEBbGs/r2bMfhz/nydPuBHDoviNBhKFqMu
gdDjgK4MrQrHsrHZ9fXU7PTnGXUZAARilN5v2WUvRIRZxIXeUGpeHtKX1hAIxSeBpFyP1RwppaEr
3IrIOz9Re9Dby0gFoyrKtC+tJ5OoZSIVn0yq2JmZDKadp3jHQjCrV8VskFUDuLfy+hswrROu9jp0
AEb/UDYG2c92EcunIb8IuQoXME3ccXV8aVfl2KBZA1W3nAteZAjoaKYJzhjGxTXO91DuCBOx3QHo
DzCR5RFbdfVnfdx209iaYun3VfXsZ3zo/3sv2BMZoNR41HERWaFiA7rjIAIcejzzmqHlDXENybf/
LKk2DwgE/VHs6Nx3d+DjumwFBYrfeLu0GvOrI+zb8saR5wm8hFQIXq9MUfRR4kQASa4TUVxUNS6m
SmzgBG142mezTze4dUIT24Nh9AMn0UQhQzo32HVlBcCK+P1lSRifZjFT0DJhRUTH4qaZvSFxzQ84
+DvkhqmWfDUWWPgRA8zfMEz5SMatBelaO/2DMp3n6sSY5MoWlfMWgUu2qfzOHNpgKOd+fKFsMC9F
PhB2una0MEALhV22qhKFQrs2Z73TbyhKaUveIyzMvkAT4Q+k1Kdv+riF6bXyWii8TZHQuH/L7DTu
3tTkt7X+4Nvqy8bPTZGzsvy8IF15U+3H+nvp+To/T7R9EqXy5CKrU8TLvlMkY8IaIJcKiYzFYozj
h7hTOUfwG8ewP2h2v/K0sVkukWZknscUT004UIifdTS3a1Z35lNQF6/lYiDIeY4WMm6Xv9siy5tf
RajfaazCa7s/h5FEMY1jWjyszwFrHh0ruJ8w2MK7oZg95v6/z8hJWs95aNmWaMupYI2apkeL43aC
mfAx+QIk72v1Xx5T92/nTsNsiVSU9Egyuv9V4jvrqf8JyLxXi3Sbf1tvAGiZ4Q3UKwG5Pc8rrCbe
OCJVIkX6nm35Y5BG0Dyf0Lww9x5U0a/Dd6tjULb2Ur+kIQot0HPa7DRTcxyLYHrITYphjmurXJr4
HmlQd5oCCHa6pBb3xYfV7H6NskcjxzW/4nXU1ctwwuMGVep9SpLB2V3kW2EX7lGNWCpsr751fDDM
3JlChyGCGBSnVL94EkCy+Qrn/FwhZM36Kk63AYZ3Adtn3HNjmxgY78Bf7MKMmOP09HiLpMyS3mpc
B6PrYEkMQA1VcWtY/KRcvoZM9Hk8ELuBGdDDhSA+18TM09+/5/OwwRSNyBXzynzJbUMmyS0AogzX
J487EjpJCFq7wOG76xYaMBzwr33WUr8iT3dyGPBjYwJBimIr4lZkgrKKwEnIYlhHlDLSWlGGS+2O
HeTk/pGV6kJspgIQ4TrSJN1u2qcO6hpbH/wJI+ShE6tu3IRGi3pZ9te/btbXUiofaifovI/XcnQV
SbXJcrw7RTgYWE2Q5AHpB9CKfGhf0Qrt4Nc3aSwB8JsWNxCRuqgQZ68i8vqD6czTnB8cPEsvFYXF
YhAnclqrXcP1c1OQmL8hz4jzLBjWNzOrlcG6ZuKdP1mC32mXXOfXucSP7oazjzlO0OInU1xW/D7V
Zf0VO+e7uXijdd0TdisDpGor4xjOU/vwA7m9N4v8+/f4iF3AS517dtImnaiUiWeLnrQsWqwFuLPF
SbWxEFD4eLo5LNVVZk8hv5c5KAW4cxlF4Vzhv/c4KAsRZMrBQNfNyAaLiTgmhgBlkazKV3rjLCGo
TxlmecFwn96wVNPlHAin4/doaqc6n/fZFVj9EKGM8qF3zvzTirDDOe4557H35iaxo+mdxRozDaOv
AEbr0v3YneNrT2kuM1U2CE/0cLMeghqZoVAzyg7Kp2srm4Hh/lkkT5jvJJlN0b7xJpgGj4y8xgD9
JDm43xtiK4jlVHPJTzcpyqLuZ8Jy6zD+94sAA0SARMMfDCU0c1Ux5YjTucbxMRDOfWCYeLTow9O6
njeOG/OGgl9URNSfDZvi2/xGARlE3gqQT2m+03vjV+TyPpCfPXuvz2IKn12ksz7mKFDS/TovAj+T
G5g4Rb0VvEcUPhPKAEqQq2+5QptCXJoLs7gcU5HGgxdRLUTYbe9GvDBgSMIkOIkwWd5ubrk0BL2o
qSjTJfnJpmKnmgR8Q+dqN8968MGa3OUu2g1pmkh7rFuoQ0RFXULjo5jmlT+eRPaHqMYtcmyXs7Gx
OaB3I6+lBsFXRIcn+fOZdj+OGEe/tAmSiL3LEdd6+dp6kwQPC84LD+T8p+F839Wbd5dO6asl3z6F
95fWsxx8UvksXZNnONKtX/Jp7lkeoozJsCrysykNTU2yoloG/cPxeTlq2nSZ6qjifRMUqqhh4+FA
reeOUdLqVAYvSR2dt4k6gdFwnbI7ztP57ZNNNH4r7s4Mg0rj1Wwuh0e67uyUd9CS25E29WAoPftD
3Ik4LJysKwGu8YuXF7p0Lm8daPByzgnJ8/bkujeE1dV3hBlyyefb7KLi318tiL7k3aJLvYk/Geg1
xq071PKvluVD+GTZ73BxJzhubHw9V1hh5/nwkNAWKetKYWcQoN9usx0SIyBr6sfo48hJt3fn76O4
oh+WuVx6pHHgGMMb33e0zCz2T2k/ebbJh/CtzLUsm7KPQlscp4YWP8xTyngAKMFt/geaQEbxJmBd
Mc7itWKebpW7/aPwGvrY/ZF6/JTSt8bRE6PrS0hdheXk0SiSseLKe0wrk/vAorYaHrIiIpPZXbrF
3m28WvBAQwd35VE2QZSIbzLV0YuolcxrK02fTsaGYJVIoTz99hpUQHmFMnTcG4nhUEhHQM5xzHoZ
WFVSP9B3s2xVOtZm6+helCxTCS6obg2ML4TRNrZnPzihjtUkhFu24nZtGXuI898+kO4b7v8sf4xI
9MQv3rlP8hk6ZljzKe6GBGh+Ik5ok+LLG0a0KsH0SESOl5gK1/4ThQqW9PTv1Nk5WVSqeYy4UqqU
tUG7bEygecsWlajoyhFwvBiaWwKOO19udb714qimciea7ad/yre+6lWYBlfhTFCL3vw2EGTwY5cu
a8NiMfxjiGZl3CNijPUI3fZuCpMZqPFV2XNNPDDBc7X0vocStIA+jMA9yswgXluX21GK177DqPu5
AEJYO59kB/ppshPqPlwWdfEjmORtnkAocrJm6I6UL1T/Hl4hQA3ewbQxriITE3AxmxJef7cmupBg
FBzd4AV/NxqjmhetnMzERGrMv//QMxdslraMPr6qPnIXd52IaFdEDebZYiZk4/yNb6rRJ7id5st2
7tP0UCc/iitnhCLX2vPdUBPL2Rn/gWB5B7LgOTH/knhm09qFD0U9tDqZEE6YAXieesUinfgNPJCT
bDJwwIx3xgtK+pqlTeRCHcwhM4PsKXtSj9IORX6pxKBMl0HX1ovOI5VwZWe0LgnpYAJGNoBi5zfb
D3pBVRljxuQMZzMxPEwTxPbQYC0O47WEGTFMouOIgFB9WNEVTI2LpFE/SEvlq0M26vO7aEjAeVO7
7IEEHXnX/NoeTVR/+kwaz+Nuuw6D8y3MgEpWj4S5ax51nXKk9nT1hiTBbRLqTqs9YoL7yGbsintu
p63cs7kAaPcwc1A3Gfu146Ti2gOln7AH9OdAQlzHh4ZXYlRYWjR9Zbq+Jeb8aOKU0b+6fGLlfY4L
uiLVASOKrJJOKssd8PDmXwJ90SIaj6Wj584wVbXXrYxWYsjWBkyXpET1A8TetHWj6D80sZZH+TS5
IMiMAN1+TOGDYg83Hg4jGbpoRBFpOPwCMo6vkAXPtDLr0Lb8JP54NxPACbtL9d7qlduHhMAK2X5k
WmVdbv6GuN5olmBySYffTw4aeX+AfVyDzFtEnAOWjs16DJHpj9kF0NCLgEYe5kieMMLgu8TIVqZJ
X5K+p3xeHfrMZ9x0xT7A3P6DJjT7yvVyU7U3nzqZbx/z76H8Jz3MX6O/taz4SvfFC7g20J7WKk8K
kSba+y/0DLOg/o97hoaH3I0ghpIBXnAJ65IiK302KJ6svMiQKqgj/K+epFayu0ZDpbDLIloK9nL9
Pjcy6GDoeKmY4ybUumJv6HQTg/WmK274SRtNQpXJkp15AZN0W3o7nK4eTO4XfPxDYPh7wC4aAu+/
MV5CjAMZ/4IcsWi0mDd9s2I6PWp5Ru6xfkZ5yhXqVCK5LvBqYklCS5oFTb2GKXpSL6RWWeLvRwWf
ObmE+83XRoPg9XDI32fehA0/4NP5FHexsi7COHlQpPBJ9fePnyMLoRdd3I6DlzgbJXUo1JNdmdsQ
mm+2nt8eEujkQzGUm0QOnmxabnWUhGtV82dvG1/IqoyTYfCbNOZq4ONNJkUlfchBWNaeoRdLCj0z
cO4irpQ8bpvZN4w9Kh7BmL+wU3NkNnO7JfaMlSiLxuKBoJUQ5WHR2g21TNpmA3iqY/H+rZCk+Wka
f85ZvMPVxd1qLJGT1TtRX67DT1I9n9qjEqmVSD9hzrwFskwinEtNerFPFi9GNaC2e6NCaikbiD9W
nN/prvgZa0NdOLLL4IaSLdwbCjmDhF3ccXSR2Sm/PHhUNmoLnnu2moJ0YsUa9vYG5dSu3leG2afe
iDX+06ktNcfgF/3B6uaQtOKXJC8xHQjexjSNJg/CGeHaWrFQCsY1urgTDwo2J8bSW57HT9hBTaYd
mhhSzPv30QUn6xlNUQEAigQ7ndxzqg9ZcNzJv9U30LiniNdv7bEq3lOd4p0X+CVraykVHJGV9CFs
aC83C5lLMA277ly7Qe1GihO+XWhw2x/E4+fNyWjBWW4bWJygf5YaWYV5k9yt2CnVHosH4l4UkCxe
apH/t7ecPauhgJQu50PpG33L2rZ+oHqojX/51K+DEAnyZTLmgwLW6jzljU7dzLUdtchRmQnta3ZI
Sqhmg/I9P+R6pJT08yL8lsrZ22mqtsgeSEn6G3LB2ezOTSYZWlqJEl3hf8V3iHpgi3XcllhVHdkx
998htj/+D4tsrHuHKNZggoxHcaIXDb8br0VPpdGytpSzHcs9d8bwMYtWFcfTiTHG8S9hzjd+P8v3
kl4ujWwgpr1C7+KviaTzIcs8PgE8HZi6PneFhaAjmwLQl+RgwqFbBeAr6vNbXkxz+zqyg5OSMHZw
qdjF+zInzlr5XLA0CNHqXPaO+XrgTjHKlEbu0vZwyOfd5p8hWWdeepwibX1wYdJOmI5wPX6q0mkr
hhDZyYPmqy1NoI9b/DCNN65CzA==
`protect end_protected
