-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
vJBAIShzznZZYmMjmLq471EYI4/bmh+AH0tqJomf8IHTkVl8LorUUoOkZqu+bXxc7uzuLRe+3BQY
jEjZXQE86etWd5C4UKdA5n+e7qWLDnIDirGi9x9cPrX2Pj5Q9cp7xaQRljT5dIoQuRM47sgFQ6x5
Q7DLd6Ucu3HrfkztXcNinQi8R7B4OPwbEns9xXi27e9Iin7K3k+6DPG+yd0n6QXsH6HnN9wO3J1k
eCCjnvZB80n/RbpTVjaUYdhlrUgzLDA7B2Wwr/4i+os4RO0qvCgni5Y8009pY6siVz227od/dUul
+Qt1RXqPJdo+0cloYHyeihjVT6AoYv1hHpkCiA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4208)
`protect data_block
2J36ITjEcHHq9+Znm3PoWzUEpgK94PDqD6ZPBRIpuotsepAP79B4IvSFWFvQ28Wgrnm4hLLzlBSQ
okjuoZKmefFt1SSWFmZz5IvHcB0bAr8OgrL8kUewOS0GsqaZ7OZJZq+GJP/6odFDItpJ3gakXRQN
8Y5dCzwfeeAxecj3gAHA97HA9Bq+CVFH7ki2kLJ23CIjieOx0ya9zedm25rn1/wh8UatdGtuOloC
uHSl/MvgoCXUtpRviyLkWZ8j+yKeilWGXriGphxugNS2hrrAL0yDndPRrvKR2uW6QHIfUwOEuXA1
rEnKI7U+jGDbXmOkHDwTbLQ1w8CkqB7A9K7/b55/Am9VQ0T9YQUf9Wmgm5DSesw8ZTvptSj7jjGI
rXnP9QFJXFDwoxSKmkO6zI0ERP2WhJH+CTsWRXk3WkYaGeunKTFq649ea7Pq6xAYU41D0d/StKae
sFXDeHbiTHgQsdLq42jFOe1svIqqU8s/QMQ7093L636VItA2j+S2XgrgSYbmOanoPqVit7Pq1qw6
QbqaZ4VKVvJJ6UGD93L1I8xs3e37OBhzOpZiZildayohbkWgVThBlhw0ghlLvJTvtAi5paFisO+H
NOGB+mUc5sO1TBGU4Kti2N4kiAtWtqhx9qJHJabxNQRhEY1QlvwoLKX9Hm9DF8+mK3yOSGpDa9vC
8ghBVs2r53neuwUrsBYs49D0VSGjTB6X4kgoWTMmPuEpbZ6MNcZUpiFR3nWRDMq0OMmS6OLXSfIQ
2YRYm4sT3iqfKzWYKySODrxHRKUnLVp2Tg0m8HnwRdb5nZbMylnjEzCjgGV3dlkE11zozSoIVeFp
342RZhhlBIouQX+pDTFXINSzIFadIPytyg9QHCkq5wVjwkbz182NJBM/NWhTWykVZUILZrxLwgQr
QJutjOJycBGw+zazyihxg5FJ46hdms/IYGw/6G5pElsJf3LvUCQsHXCs+usMMEUWrZDJr3LbmLm4
zp8EDvKyWtz6n6MHPZWZ7sg6aoyNsjfJFEA3Xohx9vIw6Empowt5GBLAx0UqwlnC0NQ3aEtk8RQJ
mClr5cXVicT9cv++WCqwkFsf3b1AG/4mhl168S2PW0DsgoNS8prA0yYBlwE1GWqtO6AezRz8qbu6
ArIzsSOp3ytZ85FhKGsVsKl6vIiPRsWFBiqDLINaQFXMDXwpZAgWEcKS/NnzPHopDQUDzooYPbJu
BsPF6Ge/7PbBGJiRtHliFhIIwt+9vOTxr/vsEbC40SLUY6Xmfth6eiyHcxELuUE5QYHzbBg/hzQL
ZIy82Wxe+Z8rdjdgh6HTYJQ4jE8/8N/AENf+qscENPv03UizDWVFdYEvuPGS8ZgI1UZ6gXcgd+3m
RTuK0lMpfBJ4xP9Aa7pgSJVIgwt7e9gcn2WCr13H065mbYmpdCtoeRlYdlvhdlvgvIKNAF0F5QOd
mMOcJbrSpFXRiV64DOy4eirKvGwFAX+Ek0FmIcJRR2R4Oe4SxF79hIpqfDe3jVjs9vdKNQg7FYZ1
0G/LwAe1dDcGPUJ7Mr1mmBMXROVAq2KMLmLVHTq79ABT1U+Pr+QWrMZ4yTy9pkPSh9dB6uiDPogO
1/uErIZmEnsO4G5PoQ03R4tRF4rchHWYbDZeDeR9Mkx5YXZxopBfw33kcBFilulx6IorvEFKc6pY
qpy3wM+tc9hPh3DAI9OmGNaQrq1yiogwMcJbDAGh+ngwI4XFUwctgzlA13d1yTg+sfv0yHXaAt3b
Zre9nxdBDsxxo1haPoPaltUcI1DpMOJfV3mHTCZqQ3SdxrwVLtyp9ZCLgkSyMYK9HS5HyPxNtjXA
Btx2NlL7Z0YZGlUVODVkTPag15GJC4yygbol2jsJmT+gD8K5Av9ch/C96gaCzLb2wJh0+f9OX7ia
935C0KD+ouAFAQhXVk1cIKx7kmvCyV+9t3bCsozZ4zGBoI5S8oJTTtfcJKAVMtmG95T/1zBht2As
4pwsUeLcCL1zJ5C/A0hR/xZI8mxemzTgfPj7Hw52YTSL2vFPHHtjYYNTjmcEBl5D7zPAByOYaLuq
0xwgYjr0nYEvxiP+wRJAvdHJXFpo6wKD+x2YmZffyL93ImIJP2U/PHaiU6fKKM/BDZjzXSe3W6c5
FnCab9Mj/3+lZUPFpemFsqtUUHoTCmyVyUofTFbXmX2TzGbjgCDuhZ2FM+2RiQx7bVd/BUCkeJQ5
a5sLcfmTWODhAQ75haz3g7uqok/yI/JCbCTutI0PMuAiCcvG1ncmP1CMtyeQRU/5JzZ3XlrQiJ+r
H91LCr7lHA76fJ52apU8oYS7CSOZnhJH+qOlop59KJ45dtutA/GAGSW+I5R6CvVlHvhSThGvUz/7
aiF8p99PxlMB0bkFgnySv1N5eZSaHxS29Tw9QSkwAxmeO2301y1ORhCQ6eEk+Uvz9CR8UXH/0Y1a
dIcms/8fDuq3BW8dHQLgZuKwdFdxZtzBL/+aN+xpPRvIkpkfox6kBNTNFUp4MxIYT6H3eVuvel/R
tOksJMbmrUHOLo3lpjY/5/YSLjdor4ArL/Xwcn+6gkJxuKUEftipbbBOqMwJe7287r9RyX5vd1Sg
W6ani/bGpjvQg/SuNBcJtEAaQLR6n1ti5yAfzmDD88oC4oCsewTERq/eATK3zuNkdqznhfLhk4js
EhHegIf5ReSvqQQhh5tXk5qcCwYvd64qsSBAK7zailJvaaMWZuiDD08VQV+8kEWxw8dTrLDsoof0
5vqvZMvKSuTm+cZhJxm9RJCyPeMerIvTwjcyyrA4HXHkhb6OmrE6E43EIgIxXA9xsH4/IZk158FU
J9Aa6nzgz9cRh4P3lveMUJiuxkkwXZ2qXfvLv6QU5k+gyBFoOwsilq5Y8rHsOJgUOJEOllOBrAdf
J7Aui0lJgVB1odU8Vhx9iMdtzn2yr5cdlZB2CSsh5PJhQWfi2tuN0dVhzfGWwNqFYmHS86CiFUhO
a+RwkEmRklBr2PHVt6VtQTfRNVKcbslAf6d4CRRNPuRy38aEg7AHbiXG+v2AprmRR+NsthWMWYXq
94PH0fEs+EkMnCL8cGV+ph/Ta9pBpZVjUQ9mYW5o9GHo1tqrTcFQ/a0HX2784hqbXE59R7EdVoMt
o6T8sqci99t4/rd5OKdEJnFOd/XBYkzqXcmvxXFmB78WajFBSPBhPw2aV+Vu2BRhLW/CEm+JIPsr
223dULi9YIkmQhD+YfiPoo0iHSpWIuq0/NZp31ptTqEFxlF+k/jLzqpzgrz9lWwcOQbo/6+03kfS
pulbGj7MXrm5s9UOFu1XcW7aVSW4zfRb1BuRL+S2IGw6I0FRo2fooX7L3bl7dynTkbXP+e8ALSq9
DhQtZmcDdoE9hRNJ+uZaNBBpUWA4vClea9LDqI2yHxycB1DqFgyKlIeLFrRIAo+Kvgg1yhxa6C8h
8G2gyMuFyR/BPwTQVOnUlNUfDeZufnPKEEMmkCdX5Scz1P3mic3EgdgSOsTYWTsgjGW9n6BcaBtV
gsgA8i9c9eIl+K/sBxBifrJqp7mWTAP6u3ptb6w3w0mUOc5FunaVjCKP6dCxMWAGo1Cx+0oOGVLW
fHrH3U5O5anIdvVtn2yQ2d/jQfSaLf1WnZNk8pqmg0/uGGES5DIILHBUC8wp/hKrEwdMoUMCdzA8
zUnpYbFySCcY/xc/WA40Oxx1f7lnzEEp+HJtJSPj9kzbiGdlka/cXtQzPo/4XxDtxT972Hql6Z7u
yjIh/hmWar/iWyPL5tnYxhzcVBnESWpuVYV5MxF0Eu0/CshW0+LTaKqVeQbwBizrmOlDxnQsRs7h
BlbtSOMG82JA/Eixmvxb3MwrBcrDN+EXZOSTRfv701W5nkCr4TNy/fYIY4EZiHn5/0utlq8GVDx/
CyQW5XzOhcgGeR406enU6aFKLIc+AXnF7W0TIPTZWNgS6bkYIYtr+4ezg0SsJn22fhhwjcQvOL/8
O/UIF0dkAnvwJsdVXSAA3WKokB71Gn3CNIZDFY5OZx0XqeQVc7hICE6nfTPNwbvOS3dNJgusj0Wv
fPWB1TnjZZ+ncD/EktLO1+7WXO+9BKH+jF6X5qVO3X1MHKamUCCqNxf325Lrg/8dgd+ECR8AiXJK
U9k7r7f9eUYIaMMRc13DTTS9p2kPfOINpH1rlwoyw8cgfCpzqu7NBj1gD+pfojAP6rrpCu2e/B3x
RV9LOfTDbPQBobWcckqRHByuS+ekgv5CNfVziJHOFYmx/HYsoD5q1Npz4qwkKYPUrlaAgHf0DBLP
Vbt3RjPtY8bIcXskweET2YefN8f+hiSE5bs2DXFwAVe+OvqzwpneLK2/65wptGDQquRFZwTbI/1g
AnACs8tf55fNRLzaZhuVjQ/JACKz481jp21fwg3nQ1UgkVBcXth3i+Knec8Mo2m70VODyQXV481r
coXYW8e+8VGQAb2lRNViOenYcIi1MWEVM/bD9jGxtRR/T4P6ERtOhmgzn9hGJysyYcIf9a3dtoLP
33XAXn1gptowfdHcauPg2YOIY7Vh+ztqq1JcAVda/BQAhKc9J42+ZZpi7Wo0qh0Jw7NLgG9S5raX
DLxHHmg41u8ldAjbhc4wfm1AO9zWnXFr3Eodl4uqOP9xz4LPl6+nt7OOHcweO2RhrAC7+C2yE/n/
1SN1PuKVEr7wWlurBC8W6mMTPam5EVh9ZzG6aY8Nx9tUWgPgA9pyaR//ZWBNCJG9sJPwWOAzx1w8
D0Uy3UpJq0wkaylzV0kY5i0lz//eML+aDK8YATr2HZrOMFnacyrbs/UanccjGVJcC0pNWT9N1R5T
suovv8hyvbBUATAdCi97UJng2b9nWVsQKWPHFCtGgNfx3tS2vjwZT1cZdULlXGWZfgxS2vJ4nTIc
RN7WkkweD1vN+gxwxHKO7k4zFUl8ioSf7tNw3iA4dqwUEX/1FrdJU7D2E95FhJkp5bG6jrVo9hnc
XvP32D5h3KPq/llI8ULfgE97ZRH4X7aP7ktJytAVBQdC3w/JhwddA9huLHfWVpG+RRcYNqduvj9B
mr2YFEHyxfdnwif2q2NXjvYED3yiwRiLtMwIdrLWBzzo6819vPzToJjkFHuOv3Bcyv4BXa1OgVB1
QxzdivzxJAQ75mfFXP/DVk3leMRfB4Ug6A2i5RsDERhO45ZiNnYbcr1T8ROk9PrHpUekSGIA+1Xv
PusGWPWYVrpVF/7QzN3cUM6Rbu0KDEY5dJryOYO30AE/xV5n5zeUm3fL2m32hfRNTcaSoA5SULT3
Tk+twpMeopO8rNuqJdxsxt18bvmncAnRL5yxUkx7oNkprfSSHv4ZzUZnZ3AwhnOKPacfTCOM/++u
fV/f4ETjgFLgn8wNnZ3TC0TEKOKbpAHJnMVReTYqUDiRsJwH2lvwgLfMmj341n8DGyQwIZCCXs3w
5dv0P6lh4FTb8vS7Eg+oLWpEJMHs+W+zjXW29fLxViRBNfwPjro1NYKyI783tJtHkrPoAgQ9+BDi
xXOOXejR5GNzpCQ2nUux31TKDGUexcXUppKYz4xpMtlNmW+82xmu9KIMi2zkWdC4gw2GblcR9B12
cHbcVKcPhnTWumyoJY2FRnlyjoDPlfM+kvOfaXWYROFWjzpYBCeu2jR8HUeShgg=
`protect end_protected
