-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
FfwaStkOumbADn+g+jXoAvjBv5Y0x8HCQPNHUeF/Xsz6fZivNmoMs3iuepoVtJ0/liWilid3KS1Y
ieoW7HcGNaET7hhEfdmbejBOQLWixF0nWgCHuR+R+KZQw42AreRSOUtKWQhTcTrNlifsDLqTxQh4
Rtn47eFnj8oOVR+Se4Iba6a9TyrSRYi0z+sHed3lvuMy2dR0VbKnU7PtMs/a1iKlmp9wwj5CkbEQ
/XbMtFm9n39UxEaqhHkqMtDtHiov5PV+FgzKksBEYGSHs2BMY/BnJ7k1QOG7TLef9K320/eakY8v
nTKSb4pR7ZXmP5yojgukc4hZ39Hhl8nAc3OHWw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 17008)
`protect data_block
8jTVfrBIbp69/jVnbMGFRPUdtp9DiQA9pv6+AkIKf3C88sjHLEtF4+le6hy9JG3bbKycMZi/8bNf
ucCAcm5pMCR9mJ3g76Ruhe2z9jcXnBSk+H43CL+TCknp9qMuCK+hK+xdmT6FhbisZe0t7JleIh7c
PG9JBegxyQHN0oKu1TMcw/EZsiGodXTYCqjEqZzWFZXS7W5uVbSJE1tEqiHkGWrklNuybu/WSBqf
hXGcWLvg7LPXHXtjrco1CLohoNg74U6KP5nSEJ0NKzrVSQ5cSfeeB1lgVE6ZtwHR5XeimucEIdpn
+Bg1P/5JI3UZS4rjawACMjLwRwjivVTMJgT2Ft/gpDj0pTFlHhmW4FlWTmGwPfMNIxSvxLqO1gIL
oxYYtFriBXU//ZMjO2Go7/dwMJ4N3giEijHsMQvLePnlm6Aw9xFF03AHikRdp6U60ECnuehDvISH
q+Lb+fuyaOmg3mY9idk2/Rcy5KeKDnyWA1iHpmf2QOgvXOzRy9YE4sdHxqXIHAWg2WbyH0XODri/
86G0EXIz/r/BKZ2VterXhehO7CS2d3AnpCKorau21RP+ab95UWrwQGYNscSdo5HZupaqvn6LpyDp
PFAUiWIoBFW7B5mi5+zrN2pxhQqeLm/IvAi3jDJkoCtLRuzoqOc2TfI2QDaoy1QUXKhaut8jingQ
2Nb/f/nFgBYzpQUXlgBm/BlWGQ6pQmI9ED+JPwG2R65HiuXqsgkGLkS4wXWysJX6tn18szHKBPEC
h0AAk/ptlTE4WWqchCO9nMT27Ehlk353/3/LqEa+8qs5t0X4Z2UvmI61gU0umjzgK7gX1QW96/T+
nSk+pWduZWHZtLyK/gT+MAf5dNGTyiBwHlX2b5dD4JPPS3ndm1xmdUH24nJbjLU3tfbW4yE9RFw0
2uQ0cv/P6++eRCE6EFKf5aCR1vGByOdteIiAgQuNcSsva4AhCxVIwlQ3u16fYCEnOujOAGeBhnPu
fZC0+AdqT2uSrAUH2qGkxtc5iI9e2tGXhitOgorg/yD7XIZvEMAa+nk4zlxFVzM5dp0E1AOBsCTx
uB/wlzRkcHxT5G9i8fchRK3IXIALKE9ryszGHwHsYuP0KtF043BmBb26zFeW0wf2OcFdWkW+UvMh
5MlQdNtsCxPkNtmKR4OBUB7Z2vwg2mQI+qKE+9cf4Igjan143wU83Y6fNeOss7vjeOx7Iw/GhzaG
UzEFtWmeWv6GjCakHDcH1xITP1RMqUctpeA1ezstG3H+1sOW3bdv+/LdmnWFWn0SpRiGyRHE1KVe
qFPV9Eyvw6d9MOCcpR+vgjtqzqwkEKRa+XikUlMz+FIB81ZI2ap+RIFDteWatAAuMrHLN0vfhM1M
2BQr8RlikfxIcPl0UQFi+UmWjRrC6BnBnr/qKrs2GO0/gWk03e4zBLR+BKvxvTVM4IMo2KpmWOZr
aWk9lzsj8quPYx8Qtxbsber1SLPLin0gTie29rNLuGcJr1yIoerCs2V8CIa3X9Hq3fW5R6nXpxQs
XYbOZFgFWE4kHwpQ/MPne7t46feLoMjDCHKP3P3Da9CRyn2EdK1EuwCBO+SNVWbPIeDeDsyRuxvE
KxM3Nt+Lin/v29r2ll4/049vHBMeykWNfcdK5PP6xjnwJ9eUws0ux7Ufx/qoCeTOMh420rcxUeEI
Kq/eOmwn6zKbkQKQN92jAfKVZP35bLvsb1Jl2dl1trmjWJBAsCvzzSlKfJIPQrbitC9SPgVjvdvp
dyad3Ga4QzJbQBoOKflsOlChVVCgiNeO6YXbpXXx8hPMN1b2151GhfEYDNMF50m7Eu4QcYmhI4qs
V/2xsIuhQXMQtun+dlWK6sqARM6PdKc7sfbccsbokZO79kF/Pf4kXFO2gUW6hFe8SQkurNzMgkBq
VfONuD8eUqgVmhcq3o+quNRYHKJOAHeQWYtFxeyheXf3/ulU0nIHWabLoBY5sPHvso0E+/E7p74k
GvLPo1dGOA+HZ/Zge0sKAZL/CKUB01W67MSh3jPLfZf6Lvgm7LjbwHPqEPF6txhJHWAZ70GbhZwJ
4gWVB03Iel3iiljgZOqDRj7BkMVytkdbMPUlXK/RYlOuNFgWBnrb42gXzfuoZeDe+p2LZbcwr/ul
S4I4v1PXIq+wSYwAF0dtxpA3Gs6/bvss3kb0Nd20SJLKUont0gMQUgFYPy6jAMO3X6+Kjo0Ec5yW
q9BfrUcmhAUKfVW6MevMCMP0j+ilarBGmQeA79eNlIKt/5YNqRYfVq9yTiBVIk5oVlWACGCZadMe
gAczMAITzNx92mPzP7Q0+fN/xwBRfnhPyXrhobaEmWqKuzvNLHiaQTXG+HjGowpSRBbJBod3qjnD
AbaUqvpZbFaLo8foclFKPuDPInoVmP6zjDecve/+iX9W9h3j4eI6Hgpign98oIAiMV2M6dt3Dno+
pvl8rcScPAlMQgJUvWZy82BkJsONFf1hfDcr8f5bMsw70LN+GgYgqSNLXyEO+biiTvc3icz4Z6gV
eJjy/ETMxElEhqkhpuRf7pbPcoS4ZZuBE049klHLOqxOTX1lZlGBdfw/JzUL6BAcL2ckxeP50+W7
qg2r9UtXUbfzR45g6PxZXOidQsaYyeni0h+pgUZT6YCOsIgi+pmkQsT+67IuePyJauT+cGzwHOIp
RUIZEytAvoK4sTKvV2AGcGUYhsLQ5eLhPBswilbh7rfVE5mje1eGk287gptwcUYQgLT+n73vEfT3
arTO0+FkwBM2Fgp/5WlVzymni/7fQLIsoLoSPgucA4bQKMm470xRi2/5pXWEZ/FGbnJuVnH32ujC
ki9Hw0KKgcgNFpYa5WXwHgobE3fBoJK00wtphESNfW+W3xxZnEuG6tSe5yBO7jiJXIx7w5U0FQK3
iLKbzblBdGObi6nPWPn0+76EsO8Pdznmp8W7HLxtFIZ7HMNvTFjLuaeD8sXnG0HVTQGRYof0zz+I
BVQnRooBltNvoKEVxFkTCZTDfy8Cy1EckW9WeIRpu2KJti/LPGyqbrXzG04NW1g4AxyDiqzsLW4Y
VuUvjtpgDaLuKrHO/a869LxRhJUdkYK14K+6dSqW/7ITKx3ANhiKo4YGjirbdgURQ/eUwWzmtyWL
Gc02EHKVx6WqYeV91pXeofb9szzFXlJKqTN6AtEiYz/S+kc6hJN3FGt6cMQy4pz4WrFQEh+7+rwL
GzB5olQ7vkUH4EpGDRCKfZ1qKQUlRi+wtJj8OivLtO3nZ848aCEVbYppKR72of/QM487R2suqr5J
cCuq7F4UvvQX+DVh2tNgEN4lhsbBKXtegKVA1Lk/+HZjxP3/WPOkSqffAZFctFZnHiOL6cuenXIW
YfgYmUvF1Mug+JkoI5MkXExWea/pWdP1+9TmNh+dEpeVBv7an0TvEGZ/rvU40SmDjLq5NGh3DqD9
ErU7bR3Gc6BfU8wn4mCPJu86JzKlW1pbmTVT0GMAtOBT/b6uwUfn4uKDIfO8EcztmSpan+MhC3+9
muTXDC4g7tbslmqBcvoQU7cLV4tvCxZQi+6IZZ+Yqyp8efWcwEiITIkOhXLmHUz7D/pMxZ1I/XwJ
Mxb8lwMQlMiQlL64Z1Cwrv3fSb/NM16upOpMNDeEh1LTvNakLZjNN/cNGs/qVarDGnpEw9rshoIA
NQF/uiX/NwH28HkQBn12/UAGDeDhpPVmauFBrqgrpFnfCZGesVwEkkrkFAoGihzf6d54PxaMB8Go
J1sCE7zau4h30SJ11OEB0OGhYdK8DVkrL00JGes7jwePq/z7Ah9Tre4OjHd+o3eI/O8UuC9GIsFq
GwKcnhpPxEcNCwGiCS0wajjNvtnGhwF/q2kNs3TpqflIFqUMqekSgWsFw3TM8ZMF5kfhmX6yilnV
qaGi26P8nxl21pVwCdEHfn8klDPHXpbw3q1NU7BpygwiBvmg4ARA+Bc6Djuza0Zns9sGvxOpc2yZ
mtvZaCoVRud2iBN8GHMrycCrlRuSM0Pv6nSOQScXJLOfE+gt3CVxWGHDGwSJTXg2YQahaKRBxDmC
KK7J3wcMugZV/rjKjimqwV5OEu/H9D2mNypeyLad+WqFWs2Dd1j6K9GbzpQR5iRmTxubw9jMZXi9
iMk4agJG8oXdT+X/vucquUtqXFA6Cfz507f/owlLUao65BfTLx5jb4qEa5+x76DMr2lyZDTIA4Wr
qHwmX9XWCjkvsDyYiJrzs3AKza+SAL1e0YZecC4MCdIAwfDbYgvEH0EObYqgLjVcfqzPaPICt78t
C+kMgx/EVnPqbDun2JWwjYqVlhBkEQImujya9dt+ZEo7lUZFQY1fRYcaZCHm8QRr54/hzmI+q2o5
PFNCku9ZlpUVqXqNMMA5v84G/jxgSRbN9chMPagSQK2q7slN8EUBpZGqwdZ5toWBsG+lyctcP45Z
pAkKZpBXnqeQgl52/y7gvxBuhZTmctJIbCPbMCeztKwUWeQYB/DA3gwEIInJfOd280yflQks7uGO
OlrIEQMhBPTqn5XeiLCWikLh1OeTuZ3EZibJj33lQgqplCuqNye2WPukSNfvy4CYlwX0ARHe9edx
X+w6quoS+gzLz6mwheeXjfiNKD5yUWoWPhS1+ySVw1Hs/j3TkkG/mVdj9c9B9cJRWgqPtS2N6l3G
0V7CH6JQvHKehWD7w0ROZr0yMULpK1yXLbcIYvmCJKzvLc6lz+hVwLlM21Wqx5nnDPiAgsn7bhsw
ISGBKIXdewgDmcuiwQG2gG3thkh0dvhpxMaAmBne2hWY6f6iVugV6yEOXL/zIfIrttErm4Uen4qS
Mqf5OxCqPcamzFdPwK3v/9zDP51OZ2wQYpKMBz+v6w8EtMhD4TpJBO62CslKy3dMSNDIEBVFA2U9
u46nJXiTJyPze41FhA0EU4EYibjuncRM+T8Ti3W+W4DYJWV7s9xTuOt0qhZsMJhmMEgV0FXQf0YJ
xG7oM1g+ZTKP7azgtnNUJj9qGPB7RfwXEiRbZ3Ntue1WQ158Dli7mp3AeEY4Z9J2vG6IxL5UU1BU
eaZuV+x9S3OTuXSrFlt5SHbg3+6Mlowevw/CYCPn++SEMjx5WRHwYqxGE7CmCB/yWXlY36/Ary/D
5gR9qJ3/JtpemOKXYxJigD6rGXt49asRRPp5sxPn44MnTjqAxy+WaqBFsnFsciU1/4OcXa1LO46M
ddMFGifxHETWY3pb7VHgzlzYaYTwOt0DedWH9wrLuodf8y1cFXpNLqYGlHCZnclgG9BokpcDzXcy
g3/GO8x6l2FWHaZv2y+hZSkn1D9n0B+ypFh7jhfxUahqbc2kGEp51WZtUeIO34DMah5DSKHoHHb8
xUGEAalBeoay1Ydszonzcj2J9slEHl4vKa1/zXSEhc8b5tCm7AhVSnRsVPVzN31Bgg+z1/tAatH7
JlgE691bkN/QL2pj/l7xEUCwo53t9jvtTmk9K7CtgrOtq3pZgGG3KkQitNfzwXEDlgkAl84f2gjR
DgE/5AqNKj3xRtaEU70x3o4l/9ZELkIZCJK/jhHpLopaS38+5WSLvZlq2bH/p0+dRZa255zoWgFW
8yNREUFePtbcTcQtAc6aMNDEXgOu12kzxoPTYi4LyK0ZNOLluYZESpRF2dfDsD7Pqon0zhQFkz2K
LCo2rN5TXNpofkKeQQWNA5GPOunze6OvANhapaPV3BU+ZQEWedUU+TOOzf2KJbE0rXH5YLWFeWp2
ZWrxT4PlJ+A9oI4AQE4G1ts9Z+I1WDyXj83sv0IUHUua52K9u0Fii5qiYVZWq9+LRIU6D1zx9TYv
p2hI3ZzrTT+gPKlKEJ5Gv0Uw6hl4qxBq6zHwRgUcwYl6sgbOSERj1TFH8XxaKhz2Gxii+sy5U0G9
OLKOk/RItyYv+l120kIY04NntNMKyWsc6P+TXVPe4xsLPqThtwcn0U4d7OqwggzEg0Bd8cwm9PFC
Yfc1bHJWE0yYuELjSu7hhF3H6K0b3txnqRt5LiONOLAT1WlW5xAagv33c/N//nhHTPOc6EAKNRgI
D4i+nT76czXE6Km2ESHPwmz9kx7ldelfOxYVZRgoaT1lHBNwANcQNHqln4IsGB1czWW/yTy8ZBpj
YsBIvQl8Y5Aro879ONXXm9ifUXMw8R7UCvGsIp3JnRJfuUg8nW5Uip9WLlhKDU4hVwMv2j9CRHyP
YzY/bMLSwhTCv3MC5cuquaxrowTuVNjk6D7JCxGhGEmwmH4kdgRaW5BlKoRy/3EZJO9FP8lF/0ZJ
m4BguglCWArc73SXpbvS2nVZw+V5tMznPmc8hiP2HSFXn0HRJEZuRxKCbvac9MSZT6CH5pSvVATb
fib91zndRwH0nCYxciyLWDZj6erIB0iiVGgVp5g8I0oqjIjE0qyPlZWIFPfNvswxW5kdXc4lk9Z2
CgAwJ27YIBOge0J/KCz7U6uubcGdBTt9uNsRLoi85dJ7RzvcH1i37oAYplPy49VM7nulbV050fTy
tYNRKKumahfQKY9Nw97tJQhiHYHtScAiLdYRum1gdptmtlA6jtJTDwDmTYUIw3+TW28iZTgLM0Jq
xqd4fbLoF9cpCfhQ11riorK7jpzQwNAkRBBl8V42k0rTTvdpyVq0zEEBUmsLXZEykn+ti/ieX1fe
fnKBaErGqiOG7v/20NsFF1ilL0PXnqOwa50L1IiJ6yCXjQ07NcsGj+/4lvvsb0ORSzlnY1hDo2m/
HtHIdJE6tQ+cxRly7CrXQVmV/PsKaZf31pLlIdHkHLHMcEVybo1DTRZzvm6sC3EuyrrTZl5bu5+n
xVqELfPqwaRR3oui1Wa3f/5K2XSB+g0rYV8W4LJiRdCEOmdm+sIp8P09wamZzl22gT8eeHl3ogon
xX+WIFu8s18WpdCr0JQiqquwqqLhoepQjNUukYflDL9fhseG+v31dK8SJR0vucbtLY821Yq8GoXm
07yYP5rKSaW149dgy+5TFlqxSPgArkOqJ7cvJlsto+k1jesxQuoe4DiV3qiHiqrpRRpMD6FXMFfu
LnwiPVN+ak1Z/kVA1CgqJDD1FqNIaT2g5omzUsjomCI8LiqFF6L+aadvJZeO7KY+Mu3C8KnHW02d
F97e4/Cj2Nbv11goyQQwzVELxktR4hHwvqF1XxAxUqpUudB/GtuIV3eYwURU3z3NikIc5oYkA2cG
fT0tbzDEqv6yd71DGbkvPj8h84pe6+uq1VYUJHL3tpE1aNgHW1N3ShElDYEGl8aH2UtJ0cO2P9eL
PN270OPNMlGElVUKeTmPRJg3tRO6GYPfDVYau9a9BdlhL/7y7F+/ucVN3QpJyrbufP2CB55TOzu1
HTKDmf85bekjsKqOYZychrg9Hxit+4Us24yPp8/3pcoFf2AS8zvROdM/oSPcrTADyg4CG93cRJ4+
5SCmpGRn/alIHpgytIweuZ8WZ4vP1Us6+scZhMI6x3fRdJfjUWaKq57S6+oohROHKBnU9ry4V3H8
ff1ld/hLtIP2ECtkt8UayMaX9Jj63JY5a6L7YbMKEEsBtHwnWC9031etl7sjDacHjgVwifaFb6Sh
qL4Q/sRpR7kUDX/0XU7RwXdFhPw8er+rq4EgC5j00FH5CO/LXWgxR3qTIiQAvn0DqzPoRD88BxHs
7E9hAia8WWdfrlUWkRopibZiOnEXCg3nsQq3TSiZSepXbLtYpo4+xj3yO2GpuLoF/XRouSqgwqCT
V5XM3/chHAE3j4qltLMCdZt18KeFZRNcfctCuq1PoXaEEy3rnF99Uk1lF3aCb7p4xmLZ9mn0E/cw
tYbYDMDR8SqXsa3atMrrncKjwQgjkmLjnUoGJWG9bsOmcWP1aVsLrvbmjaSas5whhNJpMM3k2Zgm
AhdEdTAdiH0UEjFQUwoV8HEXoY6rcXcTC10tJ/p1BU6IiY9FMWknjIj9nqdY6+D2X6NsMIbh0aTH
7f1NOxxnLUwUSBoU2BhVixrC/PJ5YMd7tTKSsNC+m+kah99ahoVamFC67q6KuahUq+BdHavWy/KX
mq88NzTF74k9Wepl+/RA/cuXFeqh3kK1ypkBBDBk9rYxhz4fpxTnAdLRcMqP78TgOJK6pup3eygf
ckLmfOn0p96wo0r9eF7nNQs2NHRVCGzoMIJF7igfmeDA/Om+7zS6OA80NdJH7jCvdIfEOj8zb2hZ
ARuyQh9Q2neXhDMdJXifC2cZdmZ5Vmed4KN/UMMUCy6dUrRabxXwYscmb/dThGhHLzinDWhsGiNp
+27ptl7cH5xFRvUR3rl++JlQm1PLlkG0Oxv5l8dxhzMJqmF3VUOssxaTQlWRuaVx/A1J3Sx/dETj
iHe36EZ2d4mHZMCj6FwPYa+73224UnTjn3zEWT3ji3BkidnYCGxjbmYdoA3lGXipyoLzAHVzLCOH
VSYf6M7/YtUTuIQ2ubWVtjxRI8cGbT7Px66YxCsyeOptWYka4yu2KP2skWSBeigqCapT5jLygt57
/wWzZxN3dUfMwpyI/Q4Bz8TcaUc+8uPtjg81TBYxSRGx8LZ8NHiP8mmZjmY4WLEh5zHjtoEYU7mi
CiUuKi41W+C2bwePTxYKI+dkwKsMNPKl7U8zFIIjJWhc/BkwOUICaSsBdVf99QukNZ9xikR29KLS
DNqcIFRsrZ71AFfh68xAWfQAtnmEXMTWqeZuTJeJGGNdRCGJPk8yKo7v6+9BpoyVYKijn2E7Uinb
UG1qkPm8C1BhU86dWJX/5UNkKt8I9h5T9k1F3vcRg0YtVXkb/NAjbGzgmu0ZB3tlmj5l2+gtGDRF
nNaFUheqNmUMoXiMQ0kitgBFNplao2Z6iIuZv/xES5WS7OPXKuLPHzLjpdEdduXREQiYJ/zd6/Vf
c4pfZersfvJscZPf8UFD1LEv8NMbuMQqcKZbym4n6uVTxcr93j/s27/ZDqXgAqoZK7VsKOPznct4
lyRQgJTWCJDseo/IZuOnfTncFidPe+/i2tK8UmvP0mwW0+ojoVhwqrzDRSBrIp+ZhFPvzenFU/6y
Es9vT3kcosKKIfmevFZIbAJ5f2z9J664ptla3jtkDq+62Ex6z/djtKUw8d2cLHAVafPxh4Emqntj
m2sHzVwhlT7Ws8JRkaLo3VSbsD805qYjFiOKKIs6mS51HRs+e4BG4VfSyGyBkjAKkS4LiC90cxcM
LluShaXT430GqfSiSSArvX3qnVXiH684BYeiV9ONepE1+p7zLFgi210tbq/vepNOo8jBSIe8QRV/
nklPZM/MbyXfTB0M4xvL9/gpg4YYcpvTdG4/02uPTtygiim07xpCylJ2TLnApwpuB+WQk3lV8mpE
a/rOlezd3mt5zw+APxjpw0kQ3Y7V7JHLWvYvAaoN94qMz6wQSAkddjfKBGjTEM6C1vszH7FA8U4U
SUtgyZjk7VesKVfgJKLunCbzBlR+R6L2CsSDf016JIoeAWjnxZ8uwYFpr5zfRwBjAOflNdxXWzPA
ECydlwndW2dknRAts/2b+FaeJtI58h2V0/bUfR4zJu7vmk1RJy8/GgBxJrFyuqA5Hfy6r6XPc7Fe
SwEdDlMJ8t/XEVEw3eE87r4v1kGa8/uMqapJuGR+DQOHFcFkp7hg4gcSSFYJNsphG+MYajVcBAAk
WJ+66PgXwcKz3XO5KSq/+kUt7f6bYoMkqHsQ5ogZ8OKOue4fGeeBuZBJKgeBChIklraINqL01uX+
Q7E15KS72OXdBSArJ9f67fdnbz8TkwshE+n99HAajpXSTatI7IISe/WxW35+467FDc4xix7wPkdX
JthWAtwZ/TtCppOORSmlF+de1hs+WFfQPQi7Iz7+TrYWXJBU5nlgbDpy7UNyda9gLgyZPMs+IM21
Ae8rJuOKALa7AHJSP5QkIvbA+JqDL4bVp2s7Dte8wKHWCibVimEb64nYcbEj9gAXFa51p+nxojtR
E+/L9FEGIyTJkYIj5DrPjE0+j9it05XjPHHKtSmFBtZpKkDyGOmjqNs93LnSQUI3ykk6uaMiuzfs
dJtsJOarmekP8eLAP5OsP6BAm4ab7qKYgWKF86dXpY6SbWorISc2eUAi6UkBqoAtbJ4glgGEb1qA
d6wquK6Xe093P5SqaZhRb+mzFs0zuGuLKbeQgVofjfpxVpRuzz37fdzykxqUyNUNu1DcixcEHVUc
9ybJf4PhU1J+N/r/VK5sXQm+/mj7egaMgQX0Xv/+cwlvDxxcyCi3FdOIVT/62K6DTkja7mdr4mPN
wcg3VNKRs3DuSvQjrvVF0h9b2vSxU0WXgjhooqLpdAH67eUeVDhDUtbqL/By/HuubOhnviyU3q1b
gZ0wIgiPn6Dt4SeFosfB2EnbxJ9B0wQwFIk3Ksa2VdMNbwBhdzvA2OldtIyv/y5zmPGTKBVsXBAn
mlnQLG40mpWRVa8t5X+cI8TtpZx7s9pOHOK2b6XFuvCf5L0g/qcey4ojFbhhjYcoFEnvdIsdMhqD
1cTM2qLryzS/BZy8wfSe6qcAHrHUCtDZcD7VhGBv8M6Cksr9eJ1jVsjfu8REH941858q5cfuIscG
F1ha+Yki3ayGdUpVz1WgO8Rye5sRiuYBzamzPyR2SNmvSAIdPcdr/VX8Td3j/lq2b9BXVGq82nA+
8ntqmm1tU3xxRzISxGFsNyIXcXVntY11aacV4wMygkm0VIFv3RReYjGGys7IudvkczRqgfeS4pWb
SI2LtIDEhQ0t2Igzhwi3M1lpoB+aC3GDOmVHf6AwUTKyhTnQ7oNfvBYNpAnaUCGd7i3Ig/Xmf15h
ER3Ok5OsyR5cMiiPtnJOFihDqHGmdEVrvNCiu0YqWvKiRrBEkjP/kcmiFGf31dLE6yiR5U1lSwzs
gR+1axFZjwFgwEhD+V+rnPRYILBAnNdBZdY024W2kz/9U+/9hndIO7yHMOizwLV6IzgBtmi663+T
j5YILxkdbmrWbTlNb7VAzdA006LKyeG3DPCu5sVrLXnONn7ACkvMwSMD3tqH2oM5RsGZx8L2aD7N
3vT3w0l+QSPkL79i7O+l8jqnIxhFW1Qz3voR6IRauIZwqKsuun2z1FAEPiPqZvGxyj0p2NkJC+4B
OXG9K5Bct06yRTAmqyJWIOnkHvUbBZbcSw88TbD5JKvgg2WS+F7BFxBLvpOldZKMPn+xVsJiO3xF
0i5wjHM2n6yA8NEhCntpH/A7uA6frQPJoZBxlrnWJVMST+KEV7siEBQOeMn6d4rzhbS9plfcNvib
lvisCFGvmyp51ghD6scyOkeaNbijRUawTo3FkhodDoH1KKT97UDRueHZCGmN8P3phN/Rt7SynUSx
kBdu0qAyO5zHKDLbE+kTEr5UO14MyQeTqG/bWo70pjv8xZh4Ca7bF2b6xevIHprZ6OHK3crTxDV3
MIMBxYGQVos9Od4gp0od/jPRQzISZirn6Lm9ZIMOe65Ah2XaLPIex0v/oRWS3c5cCVflgx4bftnM
N+qoi01o+lg3m6ZTZRjyKhz6gkTZFcO4oHzRIBWTUBciwx0TgRZXGLiBgDin/hPbx+Y6JkX4bU1/
hfcWU0T6dOCB7B1zt5LKM99yD0J5mmfulcyoM9OOai6ObI6gPJ/RFTGeF5znhz1lVKDngq+upifB
E5NWyl6Lpzd5tr0G/5h8hniS4xEC9lxRTH33AROOXbv/Fg71BYUtpKoYTWZjr8+qj/oipK+Z5fco
Tt6Yd1K4PloV5uIrV+chbtptMz1zlLamCrvTLR4m5IzpyPjfoaP7oTE4n4I6YxjyTOM29enXH9lj
BYlQI8xz6rbAEDuXtLx1VL6iPpHfuXIE0QSVTDWXI+btQSucC7tm0fzXDnrUVgboX4EI7S36DZK4
sOW7mBcqGLvcptsG7LFg/BxIHvmeRUuq9lJvrPVcIFGYL6BFi+gEK7HEf4nUfgdqda+DQaerQOoo
8gbs/xAHpq7o1/ANPSL+W+w3vG8SRBD8XOKeA3ekIvZdHhqQ1G1xCWO2CGuH1QermnhX+XAUvR20
4eHI4kcHMbzxMRX/mFbOsqUb+CnXiJO6eJjw1lR6I10rv3ZSaeS6ye7CwZq3YkE1b4N8eHQ+1gWe
/T24ZOioUVeHqu6YPvjKs/7aT53UQ12OB8/9vd0zIX/pN2yiQZCt05TqdDG3EQq4LfRKaWxZSibs
ZNJ4qPQCjp74IdZrEJelTu18AOwpT23R0po51wH32mVjbjwD5kLxN++KKL2H6cdpi4S9R/a1lvw2
Qt3kFE3GQ/3XUevRp1nWDgyVpAHZayhvPDZS/SuwmUXLhPqE3Qkvf4v9WHwz/l9Wh1EoiTyPCy73
xEqogVNk3QIBq8qWbuZklX+mYqXZ51ztSHva4S1PErwYxh/q8AieEJSyQIep9Co9lQAM58QkWvHm
6ApU/cLNOSjiBeh4VZHjK9qD1/Fqwem41l6UjKzWcVK+ZaXL0OlEVqrB0IySupFt7vnXO9009fAk
lEvFVwAoxtGpzZ9qynSFHLJeuu9Bn8cFAWyT9HgvGiGnLFVUl4XdIxr7XBmJ6dNBeiSIub4qczPm
jEPiik9YlAIvB4sV4ksEMxrdFyyLXdsUxahCXh3KYOgeHoDsAPr+DHuR2n6obcFvJC3mrU0P7rdM
fRP9pHrC8iLBU9RGe+Ts6Rd3uYcndshUsYECvwXmmzx3jHCm+Qd8vZlU+io6Tew+kL7Q1tHiml7F
fN4uNcPcX/2hrtO5laeT+sL4uowQ2ohYcrTgHGS+ifyrWxhb6eLp/XH/9uQpVqDStxILVdBQwUjk
gf//f27Yy9F4Wu/B6xtueUf+fNmtcSC4NWggiCMTz7IgWdfhdtfBNjkUTHNQc+3OdEyF78n9f7BD
+6YXISiHvFcZZjW98izfCPCTRkd7XnCNqSf7N4BI6J5fMrSgdWVGZB1QTlEkLIvz2/xgmi3dFmgQ
EfXwC9yZzlcddLusw1qWdv0VQVntazFo/oLS5lr5yv75Jhd2p5vHLbwM/QT9+yFIdvCEsQ3r6ax0
EAZeU/8AipFE6LfVM0XGPF2Jak2ALtOL/0fXf8eyH35d3lW1z/VEhGzoaYfMH2i3HipBBNGAzQES
4Hhr6n0SxZex4ZulbY6zDVp969YyqaBRse3wDedibLyozjj3VJqQEeBOa6tBtTb6rzLpjwuDX1ue
tgOxQR8hx7BATJfFWNXWRG9SGPzv0HYxRuq1Yhqx0OAgmbTDuUYIo1zirWYHYAYGPLyckOCYeFXS
DWy64+Gu4TuRMNNRQmipjcYlsEv6DBvax7wWbLhqBdrTucs0qaBfeR5iJn5lFXpFkgirCit5J9LJ
p/Udb7tiuppilJ7DGkWgzTUaOkX58ZivvTs4Dp5JdmNYGirx0qwUB0ig7HUOQwZp+NxyDaK0PY71
sszV98L3xd6SXf6R1fQBlrumVUY6Jhxk4/ThMG0Mds647aSXQmii5Ym/CvGBf77xQCXbhytGdUlS
OgfLmba08QFrroDgTdWfdVPExxxmY44M3AkMznoeag5pbeaXHH18Xqh4Um3Ac5imPSxJTtMDKkId
/M/6JauzCn0SDIZlQ1iwSxjZGoCeiqHVoGWHMVnHnuC5XTzy0rb6orpLUOvZL7g2T3+N0IyVOUfY
n21bfhPUXnkcZ3DMotxdY9kbz3bmbtbrA7BuoO6KA6JlGTsaG+Pm/8cQjQZUg6+TG1Z2oa9b3Xg0
WRJjgLHoZWxrtH1UYcELSA0vUkNysjmp5mQ8Q0zA6hlHucgXQTpTmiJf5nWLSUF4Pw7FvjWxRJwD
KVRq0Frkic5fBR3/mGECuZTPm2kwCXWgVn+HGN/FhOgA0unU+0Mt3moHdceaDpYJ1AoqV08wm2ub
zVCmkw1Ccj0GnnRgcWp7nwtlgSKtghjjogxkrCsPkDhFmhFgXx1/VNtL/GfZTdJ15uzF41erQtzQ
rf9NjSCtMka1LsTpjUlSc0JlzUChvNAY++9OKhCzoEWmG6g4mHj727QqySQkEFwzgweFP0SnN9VR
VSpyYRausImJu6i6ezJfoXJ2IfFKcTxJapK8ougrd0aWd7J9ENNjpzHcqUR051qguWMno5NNtM5i
yXsphg27L41DCha19lGUNyvDnUZUphipy60dl89IT9cyqtZXxuNosJ4A6jzx+VfTvCdEZ/IrmxYC
PFYjnNVl0Fa79KfQ8Wbi/vz3+tgczG5sxo8OwM+3QkdrPvqsbLPldNTIoMwQurNpUWxVcunLZVcx
7Mtg7M1LbAHr21LT3no9AQr6Z3Uc++kOOHkwZHAfnoIzW+HDp1FOlwuxHgwiotm6077XqsZU1SYI
Sbp3Ur70j51DWgqHJizPXQXpADjbjpz225Uk9VSg2D8EwcGO6P8OA8a9wBYWWIj8c7MZzVXn1yYK
UwcIWAEj1YJfInr/n7U28mkXcgWARLJotqnxivTv3Awp+oDXskccC/qj1bLjb7HL2jqabrdInzFQ
hzPHhi42p8qeO7loWxSIEeMVmSIrXtep6X9atexpTwUKqzmHaZUalQ6u6dUdwpUnzSUeyq67P+Cp
zNZQRNiztIn6vJHJRPlXj2Wd4MgZqKnCyeTwJParvRsrOqGTKff2dQwLsnC+6vRzkp0ZCnoDsvJX
YKoLdTA1EK19G+40vxJskFciwp74lutiiiGybyV54dCaz7kbtITGSSBdMTYEy9iu1EagwxIGwxzF
28bpDRmNMnpfLslmeWHJ9sXhJJp1ld3RfUq3heJ4e0xlW2+h3z/7VTLyaEV9272txAb+pT+ySyDZ
3yat/K42ZzGlSJBKvv+/esLaOK247JZSqkTqOk6nklRcaZkiscfS4BswJjPi2fFsTX0UetrYrSOs
kJQe/KzUE8Xrtfif5Deeor+Saiu39Xw+UrFxQXZyU6R6S5XRNyA7ZgbKzE7vkPZw9iYeOVBqrq3K
rSZ3PwWXt1Tj4U5DehjwNcWq+0Z17C5WBf6B45ZUlDZCUXwY9p/eHfQh3RMn+ICxLrPu/q3KIhOb
XZm2wDjJkO/B0kHFqvZ1Sl+H9aIrIIowkEMFdTuLgE3zHbqBhI+6b99qd+2WLXi9eEaicbhjSG0H
5GTphJgyKkpsX4zkQkbZLczAtw5NwzRk7PsAPZDa63mfipiKq9dimSU6yLriQ8NIWfuSGpduznrp
j0y3628vuGtkukQE0imbU8XDv4Y/11eZaxU5TnlaPZOtJQiULA2+fxYQCJ5UMPnHlTE+DJAodkQB
/ATFGWKtZM/QshWeodv+fUH8EZuMrD8x254apY9H95znm8FQWi+qaUxGJp/RL0wi8BB5UbaE6snq
v3532GvRQtrBwCKQYyUUwtHdJkWGDq+I4vccezteQgdVxN+kbZUMMDnDrzC6nfO9os7/e0CTP2n3
CRVxn0NrEcfg0byFOWnwVbHqrsxKvlA32pkAQ9MO4tNWKWP++E0QPtJva4M5A3qJ6dBXLr7Fuz19
FhdKF+o7qmsiBR2hmgTBHQ9wuqT1qOyv0e+jrDQJnpbU9CjuPmdLZLbD2QlUCh+T8Qg4VD3GZ1ro
Xo3x0DgdJxIBSQJ4Zj0tn//EBRpWus90J1bg5oOQa2/HbOS6XBcOJc/XcqkMLcsg9daNcFtLuaxv
gt7buRqmMXXdqYTbK46A6clHpsBJYOktphhH15VZ8fIAaZnPdKVCJ5+60wVVjVDEpI+D6fVLWd/D
+WBu4WX+QAY5CAVv6WmXZ/HMLpCtiYMVXGBA/SeZQei9Kw21AQ9ceKs6cH63zHdiniFowEFEK92C
c551RmYafOOikaRF/zqei6QdBnvUt+wmYsxESjpRcSIGw37JyrQOSoFQY3YsaQqpYyHLV042os3o
Lyx6LORcwX7ZmpjLf/r2H3DlIVqBz/mII7ZZpFRheV5Hx2xoRbCdwPDfm87u+XiphXjd/7st54RN
yzX+VRm3DK67YJbn/DenitnV4efoszhnly/8+rQkBOazy/Zp1S8h4Qf5gGde//LFK/Cdt6u79Em+
HntGOFvwG1VWHlXjLOql8Ip9I8UpVqKlhEGvO632dMxVcYQXnde+xc58TrJLpZw7/EGF8VktocSP
e9mvAWtMaq+1ghtEIui/fpaqadY4sNH4Pr86BrEB0eU4x91V/s17guoqc9/4+23GL3pLG4bFPHRh
xsdizpZBv9ttyXuxcrsXPdFneS/HfDgR8ShKTfguR7KkOoTbtoJTBnZ8YemrfUN91fliPpDab0tN
TbsFwPth7C9A2mqu5ypOJRs5W3mUu8c2JWwhHTLw8ExYSG7m2W838Z275h9vdKAEkVN4L9gICung
rEBNuXpiaqRS/+fE+4MXt7OdCtHOTFqA62VzDc+SoHrsdGLcbvLNFjCAXccHbJ5rXleYsGSU8B6A
UKC5nFWhVMIVZ8G+lV/STEKNMy7sTGoW+tWQp73A/r13p44uGdDSXoNOOum063PaantFXbXFuvHE
PPjFff+Vo1nw4vxpF35Tz0ECSC3N5Z8j03kuOc9CAtLj3RPR0yXTHH7pSgUZdRV8UTpzSDmZ0lDj
uzbH5hV63z/nQmfDuSDmHzB7HeNAiqxUn94irj3e4HvLL8zr6kX28PjS9O1jtH9Qt6u+yRtW5EsA
hoCvssPDaODhjjYvUwrZtIxP5v3jrhl5y80m22S66dP8VI4CvpBdhZpsQQsJVB1M8k95E0uuUByI
YrVZ5MMehw+MZllHUS1xt1VVqSrO4WytG3m38wIOWmk7H8SMQAe0FsqZzG/Oe3HSMCqkAgbDYu2W
g65bRMKGeXlfZFkvlIHowGYQltdNap8353asm2dmLnmvdTxHt1HMkHuzTmU5vWWP+igr/a0RYD2P
Gq0j6T06vQxhtxnpCih4Bkr0Z5kjrD8aOx9jlWZngYFky60/NQSBtq2zJ5vEK2w7Q2u5x931r7Wk
W5sFpfeJ87m0sdG3QgxvnTQAXXm8fAc6eaeQMpXkUpUmkCQuKK9ibMJcBj69TFEW9/VP2GPXoqpt
ibGB5bUqxQcKNmpKI/MKhxH9i9G82abtOrR06NnnmFR3GIKocUZxtjM+4yRmpJb96ChTDZU8kRES
uvzZNSim1hPjW21T6CM73xDcQyzsz7OFTGY7rdMLgAPPjpOrvUKhleAVThIL3fLxlYhUUXeXK7xt
UrKD3ZCc600Mlrf9r6rnKpvRfUXk8JOiEXbN5txgm6M5ZnMK/fl3X34ZuvAG3f7AKEpWYwWJXCRl
U2OGlfQa7V2bNgSSDeL4Pf1gIlZ9I4Z3oDilUxSHAfiLM81rpKKsQE+awAk47EKXx5xTN0OLgVNQ
DGl1P+PKZR8b/1Vnurs/S6KpvIbz9wCfJmVBKfNp0rkxzRLCfLCr0VbnhlljRWmq2ogi3YM0WufE
t8Or8r1AimXI6EETB4sMFKbYm1r+0RzhSd4naG2aHidZ97DFriSmQJmFTOmQAiLGkrBZ7U9rKGZC
2DARdORgUcRVEgbQGTCbplnTzUQJb4itmcJ01IpamZ733vpD43dqqe6Wb1rPZshtmn2xBROp5+xS
BxCJRLG9sIzInGJLShzjw86mRX/Bc1PzD9raMPReP8mi4oJHWKDGVBmDSWib9g+bamHoafNlPCFP
uJPWv9bK/JCmjoa+sYs1WNJYvVaFKr8cTdWHklEJgjM6zBRXkzw9pq/xkZTzoaALWW9TLDFet7eb
O0i4aQ6xWIglmcH8+uU3TyvXwqNBkR3HwNQMsjhA8478s8peRU662E8fMqzveKJtDpBgvL74orUY
CA6bkrkk88HLJohl36WTd5oBV/dQGMH5BcC3QUiOs0agI+PN5bJHT4YHxBhRa3PIqRz0P/78VnuI
p1uhwiBDj0OTjouCYeAvWfhwCXvbuIGaU3rT4nEk5kSGfh0OjnNZqC401veJyauokHRIQvQSTist
Jd5A5R6i1faDj2k5bhPyE0w1sT5JzCsf3ja8MM+xCsiJPykBI1cOtWAFAinCzGO2kivSTnGHXWrf
7bvW/Y1XWb8F5BGJuWHR89oERhIWOphjABlmXfqfuzndU5Gaw3vSsMBefacuPwPfkU4aP6rseyPA
YNEpm0SupqfWyqjeyAKKdVBq2Oi+6mJhE9c5/0+yp+GEjCpehnBYxGkbS3OXk3idXiwwyVTBt6OV
KcC9YoNIA/5co6Lrmsl43fS4/z682kBrF/Do7+KuB8KMD1hSRsW1OL/Z2ogRu9w++MHqBOU/WPZs
V6ZOjWy/63EQZSHT6JMJfQq1Jje7sP0cCJp94A9ZdbwIlsv6q/VIDJi4Avfs9/bsiv+ZatWbL4Wy
WDSHNXMno4zDdBbiunUxnvAKeAELYlrNj2KycYBvgaa7KWLnB/revMpuduTb/DgIABjkiInmT2p7
W8OVxUNb3uvzpxAS9TQuDPmv4ko7NhP90X7XzrU7r4w9AKx/g9MeEgLjGg5UeA42RIu62PGOfvSs
ZMVzwknRp7cmY2bOYBHxaE5ObbPAQ8bZj1dXks6CXNs4fwnWwvdMbgvCfhnfbiA8UKwADBXXwRGb
KG8gwfFzpRUhpMDkSGYAIfqi4NAkHr60PAt7LHAz7ryf+73iy9tc00pgyYT5dRQ5boxhqfxC+ixs
sB1Dna+W5XJ73jF9SpSMVFXqh0EjTJnrfa3hOC0rSSIauOhT7cF++16EjRIMehEwfg5oiGw0uJGU
DCd4fibW6VXvhAAc7xPLdqV+fb2gRdfdeTdh55tiqLIoH2oqavAKAfLXU8cWkKB6dAqb0a6xkdrr
nXKGYoHcmBcAeft5cXJcv/JVhvpjpwLCwgjSCO+hpvOf4sUx1oGCyihg+DOyEPNtOZANKdo3//V4
sVky0uqKAZhVqITs6LXxIc70WOkMLcK339ROCU4EjIVTJ82yKSy7Ny34PuuHSLBCTVOTY+vSOYvV
0givxkziMCVoEQrgHHdhzlVu9Hh9MDBMln5lGp+dafnDK58iRQ4at/9qD2M/VIbSRJQ9vKWzYOkR
uuMD9GeKQMXugDYwfafQjv1xNwFG4ZKWtqEvBpKSAPkHKpPIZkIFu85CkXJu110Ixr8y1z6U3BG/
QIQoehIXHD6tNbtbcSA5I3ndnNof0hq+OeWqZYlGko6tm/XKUjMaA3rRtg3bS/oSrDAeWl0CZM2V
FQFVDrYd1mXavBnh0hGAA5EERFi7b4hFESfGDJF7GJzK+nd04CSGkzpadpG5iqq7Hg0EeVRXOVQL
CpNvEP95RMd/6Dr8W3F9J8oA5w7YA4LBPU1rsrm8e0VKfuAiw051gz9Fi0LIoeP4AI90IK4vtTOO
oG/yFLJsJCsmt0tTwqyBTdQ8o9jw192PKFDOa77dBxSAT8n8Egilhrx3DWFNH8dC23vLNq6yMo7C
BYOTGGk5Duq8+e054qWf+Yq6U9wBpNM6wDE/5vZbkIo2RxgIHMl6OP4vKzOzWiVxlr2EpU9MdDnM
xcsfk+74y8sJmW98Yj/b/TRlTKePHOQLAQBo6i+9APAdyuPuMhE/fNk3jKTypZmnerFigDFNsExA
rZ5vgtMVK/y9tQT17Ub+PM04P2FHgzZWjZbKI3hiLFtnxpax6KP08Oo3egTTyt0VAVbqraktHSl7
FVicuoDyaNMW3PLbFHHT4Ub3/+75YQxkZKe82xFN2Yzs0fntQwd36zm4V+S9IcVThi6w7/tn24hO
WUDYP3N+4bpSp0OwxE0/cJBb8b9ecN+TK6Ue6y7fTc51YRgmomWq+2YRfdGQhrmi/fpw/PTyL4ws
RQ5BdKeovPrm8mQDEZfpdpB9+qntc8Bhx50vkpyRrP9/b+/pLb6hAAFBnXFuEX3W4M66XscBUAcS
by8uFWqR/AL8I4sJdZiwwX3mAAVKUiF/dTuTtEoshNX4BUVI/v8NJSfGq7z3XRK8IAfG4OJcYNFr
1bt+4Of+bOndtnla+xn2fYR0Vf1PHLGzvrGZ0PU5EXdZcwFbLkBiFTABR4kBN8vTbUzkZiiZbQ72
YOkvA70GjiNiBPTYnEpX/u7yXGVrxyckEXLt8kqEDIahOQo/VhUABsL8KRREQKk4p0EOnk/SGfms
bqKltYepwH3Qfakr2NvBSKLDziF87pV8+zwEDGy2VztJvh3RRB3RltBmbtEQoAAft5EHO7pdDCbM
Pa4G0e4xu+8jiy3ceGEdeazODejphxXvjglewpL2Bqg3rnyJM2HKXD1W2NhenGF7k5ScttZz8U+/
AmZJJ7EjMs9JeC0Y5pZIwer4+QWV78DsV2UAo9zId5HN9NzIwNe0ypSas/g5uh8RvaS2q2n7851D
9tjYKZRB8UmxTdxt9SLK3ikyqgoNzsgkcMDA24pbguye1tkhBBEmZwnvovLOuqQTEYJDrsumxp/H
oQN3GgH6jCs2bb3KyeKTTDR4ZPgK0r0SFv8fIeMyHOed9HEFgUXrVrga0cZjLyWd9r1TXz+8/uAI
jzR4xZawPrNYjZj9whPUdLITOjVMs3TWU4HQHOW17DZaDOgtiX3f7IfHmvaEOlUPrNW/Oo4KWq4D
2x5yHnqNTfai2ccoAVHlTgwqAXlScVFh4x12QSCtPGhILTdMjzVMGc5gWhHRMtk5TQGJ4bRed+sH
LC9Jx7me0z2sopqhRHbkLTaf3HOnYPjS84JAr8IDkH81xOjlzU3CUhmpi2GQpKJPzfMLflrnyjaA
VmMS0j+i6q6MFv3wQIGtTB437oHhcP9JZmYVV/Ceqp6zSD1qNv8PjHtSlnmD698yzZz/NOaLeAlt
IrNOIxyBJtZLOCf92w2+3XEEh4oxYmIwsAJ+BjbGPIiaDxm0ARsx088LSvPUFZP2H/qylOp7aMbA
nyAA5dqrPEBbk5SBQYSccbsUBWttfd0a9HvvppfAzhOJAytsHJfKxRMm6DIBHWn034L039WcAofW
FuBzgqxfl3vWzixBklvs3CbCT8o9WpdAbuBG6S5wTrapscxWdih2/OxEivaKSNqdu6Qi2FUTqllK
NvfmjJoKbILHgvmdi939J5UZIDDlrCop3PyEu9+PNEy2ZsLqij42NDbUVZRzPTikSs6tVSnv3p64
KjIk2HIzfzvXC3VXT8lexmmStK9Lxsw5Wn0RSRCMkRRfMX6457IdgFfeXvEdtsk4rSXWs7bZ2e3y
Rv6lhPJcX0z7kY2TCf+2zjKFYTMIrVxpt3BMokkGIIRuASuQxDZwZuW/q7PLNLF+FR8bDXoIwoOW
SuOZuLktgghZXrYLzS8NiQbiYQterPGExBjJXwyMauZ+AU/8Of+Ho5nOKoSZBZa6Kia5jKIErQvG
xK/klpvjFKkTFTyAtrJznQbqerufX53yel0/o88enigSqiboj3as/MGJfAG6iv+viqwAcvGi8aAr
OKclR21e1ReMZ3hJtM8RGnNQ8/nFd5drIY1bKrUkQfJvSAmomOXUjngNNpQoxEip7+3THQphbmyg
NXFkpNfllpgp7FSFUFqXMyAi0hjcu9BdDKa7sa9tObujJKT2rWw6gBxCnir3QckdEi10gy9HY1gt
yR3exolms05v9xhwKygG5wmpCKgNlHjHhdllZAHG7/52RZBGLazeOlXTEEkP6/i9guAU4bDOT3iU
H/AYluvnK3NVfqIT8vvLe+OjXodeswPyA6n3rDqfZGT7UV/+2ITF5YkB0SK1NAQeulM6KqhJMwIy
lynB9QKJvQlcC/oc0GRhWGicD+/7ffC4ay3RaI9E065/64QgBFUrYBt525AzyNQPWAAzGIzzliIY
ncm/ukmSjI7S/nsQ/rcY79Nb49jYq+pIbWQHI//bCgvy1LYsEIptWDiFUACEdM9vTdFj2OZMnvW8
qNHPc64tcjtEmUQQgGD/yt+Bqm2nNT/dDwsrikC96H7ngQRLw7poa1WYOOsV2WPs4YUUrFAeh892
GiG/Qrb31mNOQ9UDiTLCtIA31FdNHeYoPtFqIaBFbBXAD3GDEKF0Tcgh4bkTyW/xZUYzqDkm3knc
XkueFl6SkuBwqJUZE1jSckuamXwkIsacSJoteCuZ1iXMduxUltzFZUPuRtHCqkQwliN3OhFV88hj
mg8+PW8jOlHSp4wNWHkF1bfQZKUHKZouj38I6FMl7SSxVM2QhusioDwYHx4bEXlATGKXl3NcrM5n
QCmg6WaSD1EEeMqnkJNhqGPuzjR2J12kogs2wKghp6pHNPs1p3hlF+8Xbq+tw0Obx9srIxS2XtKk
GcZil9a/YM5B2ZqDNxML3+jST1dGQmcMZ1LO7LE05vjTIFn0402qb32x8cp5vlUKKsltu9auWVXX
cXOQfDB/fFL9jQpT9H+ZpHZ1Zfz8V89ILp6wiB12WfL4eMuDo3asgbCqVv0GEWN0t9uPIKhsUFx0
Elf4iCTyIfNLLH/PAxEc/hb/WmxYwzAbSx3hWe+Z03OTIpgkjQF/yN9l8QlBZI4NlsOhr6Hn/hn3
27HSg228zeg5vGYjg+t07s3oczOeWNVyBXVVmlSLZFLa88cLrE4d8phOQ4mbDbtVI3tthq6px84m
fqKKKltjQ5UQbsertxfAobdP/r2IiraDtrgwL6WbO7cOm4MLUGun/mj3lHkWVO/jcUVRQmPUG+Nm
JZjmKK9VSNVidmXKo1EEI3nSWA3wAPLmY0mFlxLod8rEyRuOHPBRxINN3UTH+CJ1Nm+9aaQpBe1Q
Odmfh6D5+9SJwIsS7bj5ngARmDk/dqq3lXHVfUSBhktUBZlbfEZ8fpZb3W3Ws6dX++PHNHWuPFka
AS39p8TTWdgC4QrCK6V2LqY3nler8QAKhQpW/M7Bk8/T1d3JPKtGjnIHqSSZI7/s2nkJBShTGHKw
T2wJpuiJOgyCTBvRzfa4w2YXrzbjaw==
`protect end_protected
