-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NtGLWoAEqDuvT2sT0s1L1Gvi2gHIMAUXIgZWO1fvQz5jQ13/6co/OAEknWtTiHUz6V9MaIc8FFaF
diWuM8vsqOO+DETg6lCPW7L8rZo8de+g2UGXDfJ26MESTY4C9d+ztsl+yV9+JEinWFZfO3RlkQpE
so/PMo1HAAAwA403TvGF/qsHm4GrFzqIfgQZw7ibcDyT19APKfatD6LN4Ogr1+lJAC1+r81r7w4I
oTNE+ZPMTrbIJBcSEFTTNExaaaJg2/O10Oa7zJYl0Ci/PvIi8YdcLfanXJNwUrM6qOr5LuaDlHAg
3/XIAf3Cr6xKVZuJCIIAH9sGcO48WB70/jbGtA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8208)
`protect data_block
GJCMPn/WYJn15PsbatXvMyjfmm54lgP64aDsKIYQ/xTj+WglYze4yHTaIQntQFyIUrzn/xRQ8fai
cyRbhWT8mM27FQrUJeyrqxNvsQz5Tq+Vy+6ise7fdg8s/gabdDk+zoEQLQ38Sv6oxhXkzy7Vkh+D
iGkiJW61Cf5ctfuu3kNeiPNfeVTzP7NMQjHVUASgztKLB6FcqGmyJ4cIDGpjv2ExSanMMWTZLlw2
ceSgMilz5K2nTlv8o0m0riQWwTGHh4sVL2az21zAyJ7AbBNQjg1xiT17TtIRxA8QFY/+iHnqJrvn
YU0rkCDCC6S0H0hwgYAvs4Y3qO1/aHgpc9774xfT4wpMhCHMI4hhGgJ+XGjoW+ZtYj7MQegtL71i
fL112xzXa37thpqm2iVx6/D5gVhJbG9FvKcb193hD/Vs1fys2MqMWLmUcqyvZl8dHfPjNKqDWPoB
s4B75P52DCuLn5Y/sWESVUy6LNhhjrdGdq4R8Q2BNhAp2ub4jXtMvfD4YnzEV7mI1o2+1elqvZ8E
6KXkitzHs/54hgPv7LVEbDjucWyn/dir+xhrtilC7sWtdbXPokpMSIeD9p8bySGQ+x1Los+nyGcq
IeAlUJVcnxZTnEl6N3si8BztclzZNk5nYv69gazKbmAvhS4YQvKXUn+7V5bJwnNQEZGpZNoadQHd
AeK1DcH1aBlgJ27fDxiqiPLFOeB3EwKexWrcIPCti+XXCGXCG9KZ/s91QDp5Mifc1lqKt0WWX49r
95151/zpueq5vYKThedS8S0ieuLwDsx8UsprqzVqgkhvzWxC4RAshPA9cLOo+58dYXout77lEZxB
/m9LNKmjjt5DuoTP2AIPGDXGfxySUaeHvDG9kGgFsAwxBKMF653R1DKgmR0Khbc1bbSQWfOZ8txh
iyyg4g/30SZg3jCVQCyN0fuWuEHvkIo8yfPKCvl6O9oSvvh0A7o7w6fjc3xS1VWJIiH1h+U1gQi1
sVcO/5IKLcFvRInfFSRY9XxIEep+1ivQOzQaT2kpAilhoKToxNEnnTSwvxcnYeJS9HIMuM8ZFEAN
9hqDDAh4+qWIi6MLB4IBwFqkmipAUs7gUgoQaZFYoQAlfems3cQZfdsSNLxruxkR4UY/ca9KP6GK
NGjXGKNwhji73kI+oRi/kdBF19fcD7uno174Ja7AQunY+93zs8muEm0bLyXShT49IeeWAnGNWg33
iQx/QHRPRKdzJoiZBaRzKsN9ZyEKPO2b/hzPlmF82bNtw3cuZo3/ZUTntdxMeC9zy72qt/IT7086
kqh5MC5wkzVxLBjnLCfyVTZi6c9svX7AVEeayg5Madjxk8gRX5YXJdq4K2QhvVPGiWLaonr1fyCm
jlZzfyfTXpfniQHd4vSWRXj707H82xaF4JQ7zL/udj2Yhgl2gblKDOYRSw4NpItdqp6FPiiZfIpX
YlLA0YK/X2/XZqWORfQFNVGPYNu+s4TOm6Q9qQtf5AQ3coDABSXJwL2/G+T0K3wFQT2Aa6ItKMUG
XlF4AFWoEhXQHCNBcDT3vKYWQmN53Q3iNt3Jz5MRf7jSj4myOM6n7ODpgb8tlGVLPWvVy3Bv/hFk
7ap6YaFADldeeIW5r10ufHcGc02SG1UlMbFW6vYAQq8K2N1ERmi8jCqf2AGvGXhrHOhN9JM8Wt4J
lNNi9IOyl//vi83+IY+C844L+bNO4Wr6k4RiE4EcF/EfJ1rQ66WikytilDCDyy/NxB9BXo74vwJO
sermnAv/mAsctwGhzZWimfviN0/HGWZnyLb9E5HfFppx1WV2IB4UbLQF+P1gPnGYAsWpxajHsrns
cUPm7oaT8nznpzFSDTbddY6HSidxTstNENJOUYZwlPpKpnPRGoB6O0UD4isLr7/W8QCp1z0/30+1
s+UlF7W5pZ75dYwyXnqNOncmU8cfEs7mpFhELquVi1qAs9rO3CV1RW2wwVdBsjCP6QT7FvE0Ej1F
GZj6AImjmbbmLieFebWW7qid10byvyYKC0PfX/M7YfV9TyUhjj5LzNAZo3v+5Gt554BKFLb8eJiG
zArzScmR/1uDBdVwduXI+idIomi7xUdA5b5xkEmAK28eNczIvzLmKNwrt9uOzjLRvjMriymRwzfG
tPECbDD6RNA+yFgTHP57vb3r7xJs00XwYSiwmvOpVR4e2kkIfI1ItrB2T8vw/5qbPDWsmljgbjvq
wSEES593v+8bM61yUkxEW25CFFR/24yfnJ2dMQOLbbgmPbTR2VVriZ4G97scJ/7LS0dY0ezMltTb
YYI1wEenq1Xn7qrdCmGf8e8zZh1E9p4BbXSCaWtEz5ja6NyS9AlyK8bMx+whSnUHh0qsnfCct2c1
tVWL0MnlBCtC7n5ybkdLyRF0byRMU+zfT5TfXPgTvFkDeQwo4WFEdupfIVEDMqtAFLEUHJuFmT5i
skWrWh73bluBKNOfIBseUUK8i3cl+jv+2jag+CgZKpZN8CglnYJGeAPWHXlcdN4yY2HMChYsHCOj
mFIjT3nQQFn2kkSGtAydUY5mTVBg6KrkWZQ41eS/ydhOGRbqp9eDZ5JDVO3DhAcSDaJ3F9xDRXC2
7JluCF+yhhjwPC5936EOg2DkbYI+FKSrCCbgJG4we2HO5hiIQUfCq1J3ycOCmXSB/wix4tU3AyTX
tNZCdvX96Nv4bW3d5Exxm2Ch8j9xVF69bov52tlEkJWeYeMaLqLoPYx7wCLBmXFwqoC1p9EEOFDO
omo0+Y78LdxIGqWP007tj7ThkNSe9tIg6nVLdYuFpy34QqLSAE8tPR7EAtvSk7YbgnGnyTheVpos
GDz4E/Xj1isg96BLZ2FCplPx8hyK2OtUoXSyyhMene/CY4wt8ll0/X8e0JDQ5d7N7Qsi1+A21o5t
nUynSA24PQheA1vVC+yInS2UfHMIGQal60ALdfVKI5yt5uLBaIdWa8zjfARRLooXpmOvz6elokFz
py1lhzFsQB+Pb65i5QnwDYpdofNLIYXKG3ghygFfr7VfPmzq/qQcojrTUPAcDCSGPT+H9VQMjf1F
9M2AZR/rFjTZ8LSWWnmdL+gNF9s8TZ0rAB4hh9+DuloUSSbba9yeFebLl65Z47Zel43BD6RyqbuP
KrqhiCyzkcuzILbSRjKBlgC8Y6XilARUd8vRe0J9cnWqGBStBCqbzD0TFNV61sDlKHRxodQOIv1v
nrguUl6P4LcNfxZb9P6pD+QckvQCcXV0c+exgPFLmvz1FmB/a9Ez3w/pmlBoXfi6816x0GRsKljX
k7ANt24JX4ngpJbVXyTBPMB5SAJacjQhsrIREF7p4uoNpmtUNsb+peAJFSSgX7oSulRdWU2nAzad
rEwMZsPLTKnVPcpYUVmrSsf1vK8khWjX+5GgQnPIar8xIN6ApEft5y01DpqAxzhybxilupIO4r58
aqcTipk3sLO74bycEK+ViyJ+2B4EgPDfbFnxX3A8UWlnI5cpkmY/QoiA7nzbaIsr6vnNhGchi4zF
Sn1YJEjY/M4pmmqRQSgPyra2wV5GbdWPgUjtcFPOcihAnqqTUfilxLh2ZVPtv58KiKL1A3Vh1Grb
BNin9Cnf/G7Iuk+aohYjQ5/95ML60HlJcHo5la1IzhXAp7ujvkaD8OYxEBtOhdo4ZzUuG8bTApm8
Sy+omL40zIPxXNXkTaMjzZqvYe33BJOh/Lyr6FOgQNs7ThSJQVTJ3TLlqNM3wea1zOKOv2o/56HJ
qFxp/CsB+KIVe+mjvnGEoJTpSU+cmQed9VHiP0nz6P8YRBYTG+MlVv90Ae1UqcqS2cy+q5iP1hXl
rFn7C8NSQWcA47X37+PlWEsE+zRp0LxOF44/6uTCYyOsybv9SOQoOr4OfKa65dM1pwHfURFmfHAN
L9PehKUUKpvtPTD7shCS50B5//foRriOaaH7h9xQNXpm6/WqBzrivYozLrR4OkLnrPTMONaaKZVd
d1OK4epXjdD8cnc/+CJdsCJIWUPdQUq6qvKPfTAbSwOxADsl6Edg8SX220BYLOYjhvNcqwawmRnd
8qQdHmplOaH+KK4E7ukNVZ9R+UyAoPM+dp5LG/NmYfVlzMS3mKBUea3Y2HT7/sFB0JX3fsfVEKQe
YrVNY9A5sqMdOwIklVPLIGW4zv4QoEdU+mtWm5Xw1SN4luj5ayOUwhL3jCjFJXQWuYzS52ERbwp9
+KiPaYhYW5hVoyclpnK7oZg4atb4oZ6ZWooS3XUn5wHcnF51S3304AAPIcmXi761VL548WnTxrsV
EusXIBdOHWaUW+wZwuvyPX0fsBvm87K+YeAVXGPE5GgWE1lpefOwXmSezPKTyIv0zdr0VhTE9DUW
2n8PIS1q09afJfpymLxW6AM2SvndRK8Kix6c8ew44IrH/a/inK0GurKYJz07EOtpoJ1eqVs6/U/H
FWs8/4HuM3KJ/eYSjmNM2Wq6AFWt22YnfAq+WyzEqyoa6/SgnoSMiPv0LvyPoDYEHT8otWazbp1u
NhVz45cvwbOx+DdBROZYSvEdq2/Z1KPzj/lpPnKZGBBO9gb+ewpRprvLYiaZS1enRm36eNENMoLM
uD5lvH6yTwAl8vZYrI8XA3XEURkd1omWOiNLogEYhgic/iZ/g1wXr3oHJftipoISnvk/ofNLpx4+
KwuVaB4ifpJKlbaXyrkDEcr9INiYxrL4ZcpsNcZksYFaX8rwn5anebQvpou8xQYFhBbRwZapXB9d
WFM+iueB3HBQkH7i8zhKZCRZfANCLPLb+hYUKOxsv0J6gBYtQOpREN+nF0+r6zYD1oMZMSctH8nP
a2Co+h0dSOBU6b/o4aSVjaRs0PPrJvUL9NppsvB0Ut5luW5cPVW24vc0T4b2Bnm+KfebhXjxJl81
CqsS5G89zOiTBOTL3lvataUT0QmnJF6rrVfVJxL6bL4ncZa5Krw39fNbrrI014QlbbXOd6EK/aMS
7J9fGrUX4FPgymtTVv8PdgRqvYit1VONtiVvKAkfhGtCyyk+fXXV6SnJ1q7vAcJAyNtsmZEvHuau
EpacdrNCC3AbVz2J6QWJe/OEZISZo0LXf4bZFp8YqZsCxDg33sf8xC37hLyeuVO+7F+hQztmGDX2
J9lZdW/AGlPD+J69Upj+CTubIRPLZNwJW+Ds3pFuTlcKQ7U2weT0DkWtddTi4LS+vOf6AkOGRKnR
vws4OvRpDjZWFRlPSViJybh0EZiP5+/3ylnuNZvErOPGx4uGBplCk+xLIT2aeL3E7hMnl4vq/xJy
/GI0sk6N7HRB0djfartC0rSLEC3KXmJiPHFMmCJ3KbSJ5lmJeN07wEZw0rYhDBRdbkKmwnXT3w2N
VMkBgIwLMHgIM9mj5PeyYL0iYNpFE7nAG1HD2AdSOwYyAUGNnPUS6pjDCnl7ctZARI5odNG+1gIu
cySb53bw35oT2fxENPxuPMYQRjWv5zJqD9houekfiV8NMJRgafGOelh4D5qZeNdmOtj5ugK3tCgC
HoQo+tcXJMrtldrDebikKsZHligk3Gail9RolHIGFddL8LdwAWwbfOYFEYpzJmqTFFSedX0EzHCg
iwLwYLW9lxQKtAW/hRRWzQ+iVsVlLEJlqoN3rU+Z+lzQoo7Brs3vKLDa3EY1T4OtMIc1YojA7oK9
1PGoJ3NOWBEI3fENmFiEsytMCuqGFjWeu4imSDigKXAKLRCdVaw0GJumSl8zyXzA4wE1/Hg79/ug
E+CdbnQ3TSKjyJi6ug0ZNtDeNmr+dIyfEnnhEJsPabS9Gqv/wVx4ul2V32Poo55QAybjlNlnuc/2
qgajHtcBqhrHTTtJvKzJsYG3B+ZwOhoSTAE3NAHUtEpVW+anvNmsoGv0Dyk+3gEORtVaK84SNhYZ
lZh0IcBBD8MzaPKjC8t3lXgIf2NvtiC0MePcPJ5uHv+aasFlexWEFO5U4403BpC5fk7QsdKMuPJK
hZpiJlNDUFEX1wNVM2PjM14w4//2RtFaMwODr97fl8HWvjza+ARLMSX/yfd3dCi2ziycglnlHBUu
lBmc0yjTBX3ZYYQzg5PUImD+4H2grqTzLrhIADbHCuqWspUfqCGNw0DiZIghUCl2TgcVp22MQmQd
9THms4p85+TQSnqq1rJNUs6AKhbqP2Pzn92x8r190wMizE+w63Jr4phbWt8cDTWnjE/9e0w4QYWW
97N3TWGg7UWNsrNziZQyD2Rwvrn5q/0d1VGnPNF4j0bVPoVHbw5eAwgtsQojj/vCMkfQ1q097a4R
+jU+nPmyD0ORet+nc5CWfCiT81YY3qejjlkJlwapn9enTiKxw2+1RQ+oxaheNGYRVujadIklf/TT
wPD3+hsQh8fEXlLUmHss5HOJQH1H8Fd6FWkMJMcYWNLIkfnr9jKRqVncMUVWqo80Rqhy5mApZavZ
jOBxgOMhST+sUMc9+g3ch+U4zHdfXgJ947WEi5o4iJt6lEK0HO/qDHIBOBEyUDCCixiLQJ5XuVdD
eP9ZgkeApCeJeaBbuK1XLeQJRp0QSRBbvmB4KjbGIh3gcQAaEYSXnwTCqA8CDWdSIdkJMzByI0qf
/U6/yNHbeLINPr19c8wWeHX/Q+UOb2N1KVKoE/OoN1y6z5hRM68qMcP53cqjuYP8FZMnMcA9r/Hp
RN8Oq2/wep7WRdxfsj5z68oxWHSDN5rMcCkzj0ymCRiiLxIouqnu4+w2gToKIyvRA9Bj/t4R2H4l
KoKXAfakMg3wUQwO4DvqYWLGeSROWJFapiwrHCunxSYd70rKDew89eyao9qhcJgg2bjp/suo2S9r
vKe0pA2E4/4cwU5KrIXc+gPHz05+IxoEcnYzmDhV/92a+PQGka7nXHUQ7TN4mApjbTHG8Icp1A+A
+58kSxSnyYs5+dAYscPMsTTSXbj3LCphDMYH1wF5Olpkq5WErHvKj5tk2oPFbISVfCJPZov9JPRb
eh1IDqTAc1lf8hm2CnFlgtA+9NFvcU2faWoreOLrhPsy86BhdRKlYWcr+a3OSVucS5XhixY2mMQL
32XJ66lwqMhTxRu5NPhz3Q/sCfo83v/CF16ItioBNKOygc+ahItA1fxcQdYNK4COkWvKwRlcnLWC
hKjcf7laiAUuKguCLmX2NPwtypRyuErxcOQ/P0DHUll4P8Y295gu3lu5tfusnChwcotmHHjibSnE
tRtO/PdjspfwBWq02JByc40VoanOa2z6peBRxFJCfyT6DljKFGTPNL7kx+eGhNMROjhhFMYv+236
wtcu0QBjAsj81yX67nUa88bWL1XF70JgehgVtcnD+esfdfUi7e3gtoMsrXvjmeaog0fv6+PZsGLR
R8KN1DHu6zk9Sy9FRLUXm4aMYrb04M1299tqp2Gn4erZp6EwUIS/0/RHplpzzx7hneaOrr32m7TG
9Ppyf5yggMw3R8NDnoAENyyQZYvVdh6Ctjerw+v0UdOazL6Evmo/7F/ifEQAGrS+S4SJUq7YxPyj
pq+QphYVdPDR2ahlHYcmBYaZalLvuaAXjEvl2UlNFQT68BlVYVwRh2JS5c8iRk09S68/t0jZ1rCX
bnCpXrEqxcyC2fv2Wm4XrjGJZoNOaVEieaVZSGE8+ql8qlemHLjy2Ld++4034Vrl8jFcdfHTTOgg
ULCEghEb73lo7R+yIZPGQ3Z0kxbEUUonDDXJSx6KeOFyX3QojeUiipy98pEcKgs4ZlqwWUtl5Lew
19Sc1VHRPI0QckC9SIuRksjsZVTIxPbtmAhi1CpbBzSnzvxoZJjGaDKdldS/NLZ64niYEv1X+0bg
lr2kOnrMDN31Tmfc+kZPgZe0k0JtVs7BK4e4usziYJ2qvweahDglGk8OvzLJ/z2rinIhO8DQz85M
bFEXQiDm7Qd8TYr8wRhz3pN3TxdiP75wOEXgjyoHM5EXvCuUeyNBynuVMFD3tmAHtwngQ8zVgXOU
ajwUM2l6PPSVcYKGi9unrfQdMgR1H9vOzpJ6CXW263sl0cWHT5MrWlziJ7ctI+9+XAnZYCbl6Qe/
j0/aNxMHBgxYbrRBcqsHD8zUmlFRyghxqtnvuG+UtfexUbyPlXCIZ9vi15bI/f32mdTQ2Fasb8gj
ahJUkNl9BMt4BBvSuXhfPY6x+u4ynVnHOR8m4MWGjgwA1oj6RmW7jF2anQvy3+q6xpKwSz6qffhJ
JL85fH35/pXQgQNi7lOeaCvPVMqF+ybQNBzV8u8/qUj5fpgJpvH66UJb5+i7IrXogZvfSHguhqdy
GqkEBKz9G9x29wpMCNppOIRu8nX0bvieZKKrpmV/Q9mCus8AWVINziilO7SMEUjcvZYX2EDbdW2I
0OTYp5gTjs57hniWQ0knPAHOJvpph59B+XsJBcFSyre5SXK3JKvRj6fnzl3FY7F3OUkY3fXqnG/y
+DVi3HEbE3PKIJYqMwvpS0DV4lao35cr3+h9jcav+cdZ/G6Wj0njT1SffG2VAbAmTAQhJEJI48al
HnAM71sqvHbXphN//6lVQQqlUAlVcfKBSOdpT6SYG9Y/uaQCht18BvgzAUJpchjK99GbEY9NshxA
Z8xx6+kC18IKBrQEllJaalXXhPVLOMFHFJ0fjy7ZnV1wOqUBOPFPyeXUcyjO4DApy4isdQ7LxbN1
Ncq7fdT4KibyovwqdyNMPa1eosgcSAs2rw0oKYAsegkpuQeGk/hd7G2TopCKZ60CWuJFESc6d3MD
ObbJyNa8I3wjmkc26pWYUG9R9cwbm/SZHQT/bFAnumNPtCvHLgPbXE5ghCVcxkJnjwpI3S3gaNgn
isrViTAGdu7ytW9XkOqIaWkjYAt9H+YoYW3xt02Zu//dobAOXr0NbYJ+HnTRc02s51QTAeYeGo41
BrUT2gjiTFvyOY7jeSZd3byIxjHAUpB28HKILClqyBCZLBQwLUE0FSK4E2sZD6q8TvhvJE7eR7Yl
5MR1hJ4FByDFJZ6HIhcOiDl+8u+IlLwgC3jlibMVmkjbpSqcsK/Xm/Hj41jl0PqtwsdMyPHVSf+r
0xO2ykGeoTKYDD0H7Sm8G5rrrvM0egvSeN/k5tWmd0FKyVrpqba6eDX06eSdJBBJmXJTPnStjDOg
PWX3r1xU+VXPvkcOJqGNZF3NN81VxvKNQeuc6QXh2i9D6odjpHBipgEw481+Vczp0DJBaUmnrvFv
0X6lFVTs8Lx/O0TE6a7yi/v9Mvndhkf7ZJuldVGoKsX4JQaN44t6vKaTiWTnC2E+MuwlHS9oF4L7
QSCl5P309nLq+IffbhakkPlZpfBd0NDeDia7HGfqJzzUW5adPnjyXrlHoV1OgBsnrrsRVkPQMFzF
WrBhrQOjWPWuxgru0BmI9mspeeC8mfFg7gaEZEqgzxhMqyUF1zUC0ivNTBXgx1z9H5e2mq/BoVPz
kaEkWovjKHLECDNC+gJGb3jZyDOHaNphInkaP6/zAgo3oPA6qgVrovf3s9Ue4xcyIZPMROioyTuY
au+lZc7n4b/ZkktLgR0rlfUxO85keyUbJSFVM0d0QN/104Q0/iG8uh2I8lgH2dkUogPG7yfcbUQg
LE5VHxkNZqPiPEpUK2TfRFqN1fdOz/l/VwlyDpvvkWTZFMZDaduw9bePOOIS9uqJMNL7mPx+dhq2
QE8i4lsxjViZlJ/QwIvo0iu+jEHkdfIVu2dVL9O2nE3YZTvTf6bS/nVUt2IVGGYj6hBfaHNyIQEL
n1WRImfOhGlitqNISWX2BkhhWRXC9sJs2Qmw555LiMfnWBNHsUNm/W04gCGs8Pyb5pP8xg8XHikG
nRSELtR4XTMZ3YkGvXGxgvCJJOxRc+c4plhES1zHU+7vXOPG++uENZ13kKF1iugnb4uBbhKSsbFZ
tmgIJN53fkcAUTBxq26oolc2NvotK/8COc2vVhohc+5Qpw6+I69L1Wss4JEtv0dKw4ZuT/2Q8FiE
9prp8CJ5M9K0/FohAlVkEY9CO1KEBJzIa3BYsGLW52h51ou9vJkj6S9c3qoBGy7749BmXFVcfgcr
6aTyU8737myObZfT8L1Gf/Ubvms8VTdAz0czaB4GpZG2NQPa7wb7lu8n+BGFZNj3PvYXXWHsy+mo
EbhGTZoo4oJBxVpIEk4P68hbH+3biScoFVoJ+3481yHvvteLt1Oedt4RZkrHWZcQlVd4MxTxLbWk
Wx8impkZyWcSyHPtHrvYXlTOzei0BwdOMTGzk/dJUXubFIwSnLGFO+amUo4+dql9kJcAgVS+uvV5
TmaqvYbEiGuSl+PIF9bSrlQe00EiAb0I298jVC090h2U2CyHjSKvG6ukPyOK/xsbNu3mgSO2pHJ0
CjKiT83RvLcqz8c12AcdxrSWt1MiBYL/DtWdRtCdHGuSE6GHPu8pTSrbNedCW9a8KrifI2MZu+NQ
Cl6bhoK1M5GXDWuU3Miu2xYwbGE4dxDITG8pKPV/OET2goltUUNHePMX/rbrAs4UTEiu/RCizbnj
IsLylkQXWHp7IcAmC4UdPS5D3/flvn+dk8vASfFJTtP5vx0QCnbyn2uNix6p+P3G/mY6eNRUVpXJ
ewddqrMWnU18bneViSvCOOL7k/cjRObEc0sRTrfV3sfbIipYfYCFuSLcmqSMsbo9AribRkb3aeK7
i25iZY4ijQNp8SdghsQ2wZgyLnRBq1rpsgJIBS3qn3zlsmQa8m5ElxT/AnfH+ZQrTmOvE+xjASsG
ve7RQItlsSN6X/QMqPZeroO1yEodGC1w3nC68IRHNb6tcqlEIA8WJ2cdhNIq1wSELSHkuUFyDgWH
7pTU04jzgt1UFM+l7uRVRX6iX5Ol+aDKbST+fMFfFznOwH1H8XnWRzAS5ekd7jC6KTxlJ+vDOH1m
hdW+x6F3noPwEsIRAY9lzG4Hpjlj8E6N290Dg5edy2F5j/ArUMwRPwtFx6QZ3G2B9XmZ0Z3jocuf
2EhrvnqNhetZtur9gAt/OHjaBszvhYQV7/GGHJU4h9FjSxx3Pa3KE+en3pUVu8iPjap0CAtPCGSt
`protect end_protected
