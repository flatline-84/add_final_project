-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
GMSvSnXXYIE/8I8rWQG29wrQOKKWLTzoHlrcbydP04BFlprBtZItOn8M+KNh69XVk+wkSD4Rwx9j
7JGU4fE3/Mo9Kub4iRNm+56athVPcLWPRZjxGQmK8lnxE6vHFFq37Bsm8omf6vl5oeQ49pWna7b0
SkD7p1SBRPNCMXu8g2NNzuhdz+/SQTnf+CBuP1wtdnEvYNG9V4UbNDDSDxYxY/5H3xBycHcGrREZ
sODd35WzT5CouROVyBYrCEHY/g3HA8iNLCoYKzwwtgzuh8uVMGCioHzqPhD0vhPe6w/W4NoENzGf
B2kDi9J77kWTsqskPNU+ez0NqR/9KuEFnkFJug==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35616)
`protect data_block
Qqei5X5rChXUizIOZU8CqpYa7ooWOM+fmDiyVnN9/jNo4k9vEhlizmqYZOctIAOHJD7/zX94g/HO
/MnwlPn0ERHFU0uGakXY/9N3GcmE4ee+6BdBcGTI1slCGigu8HqDnu2dkgMJGe+iy0dNiKHoNAgP
LGl0nTjdbxr1IK4910YwKja+GgCqyfEpwsjBMAGl/S4p4F8eOYJ9yKCLfeKN5d0Azl0D+S4OTCiD
lJUVF4A+5b6wtZWE8z/TBdluFqLj/gDGpEDUQuKC7oCmLS0N2Hwe6sUA6rgLEms20ma+GmR/vAZl
HX2tgJ0yqqH6zY3i0zsO20HuW/mQ9UcuBbyY9tcV+G1KI8rXCsMH3FqFyTYaIWN8hHDMPrv/w08e
LD0rjV3I9DYfxW89bdwPVkkGIskQszEA1Bl7qXbYCe40gXsAOIjHmIuPNX9FdExLS6vXIQ4fBqBG
BCRorrFy0FBg+pIR6CYOTbI45HmVb3wHFD4+KF2KEJWf5ZmuzgFyMyqw4WKGqENkkfDoIFtgk5bq
QWmp7PDC7BhAzjaQ99l1S/d7sXma+qKkIlwtoPpDM2J+mZq6OAj/mpz4biMTFmh55YtvIWOL15m8
462fs9Us2gWlkwgc7KrnIgfFhBlDMntm6XC65Q3wzcz0RiRPuqhf7vyDEfz8dB1qVlBG3Tu0w+r1
CIlBnEpQgnmTHdCe5SotuNzDWp3lU6MX1hWasp0vha1zmitWGruZ/p5+q1EST7DNPjI5eH50hdK3
XyCOcxAXEOJCtx7PGFW40SO0ZrIyu9RSvYPtEDanO+uAlzzS1pWmRtS57mMsahGoUV0bDEmJB4Cf
IXR5QkaA4Lx9WulhRFzmbhONFUmOWoDY8Adtd/+efZwNRcBZNySwgCQziZ721VXH5VbPIjFAMYSD
iEm3vUv/60F0Q2a1TEzwYis9nG9GQrY70yrYTQ9eBagREuV0p9CIQ/qdId1hc7t4cFWVbYS3VfoT
7bCkGG2FqDajuNYvJfDFY5H0U6RKG2wkca+6ZrV5pvKZOq0lhJ4S4Q6gc5nD4R2bdcO8gojYAn1/
pwFnLt2MxyHZZ+fhtX1ubd6MxIoaJS5I6gTFFjMvuOZAKIOUuQGOQ0kiLLZzYnb2nreUSQjanW6V
my3kdcIB8AirgzLUfjpaSZnpycpydZdqc+L/GYdz2XXko/1p93TbI6ULI6XiFD2bfaSEwdGBuuXT
D/kVHyPZMomOtXuWlyLt3C1XRi5tkXeL2cns2kEYv2D6cFH3HEX/DVWrjf3hypglCoSiSO+KJPYF
QK+1+AQl//QwQW4nXXqqHFB38gM3jqmA+KPURdx4DD5ZiBOrugezn7a0drMwFjCrrkoRUUq1wWRi
LLnTD6hMUI0ETZKLMPJhx2vN5jXerNLjN6HFKMEp/SWablEhzyUgoAT3JAbVZ0j0XoCNKiqxpQxj
7Wg2NhzBsWec2XrHlMnnhMR6v/KGvuR+j+f+R+akYSbrvEFHyZgaB3KTA7TUSusWMZjFrEpo8QuS
eyf4qhgaMY+ubYE28tCflj8vNCw/V+TsanMcyhRZTTYxEfEL/iOtrSJnZPNyZ8s00eFs+hXu4O5Q
hvhpGoAz2GF/AJCZgMac3+L/2RcAPF/A3kfaeh1etBZckf+2fhFHPxTi/2kePLp3sNezROyd0Zdg
lmqa0pmUCkVpeLVmPdxzoeIWgAmXR94P9JIYJ5/6gOrTB3p751havct0SCrh9Y0nV7/nvTYNJDH6
7feMxzEblE8SuYI5iqzqp07pmGXHDhdEyJX+4IVuDdIbRSD0sG1y8gXPEzmSeKrksiNcItsBrTek
EmyjQedZ51ElzJempYQNqMKYzsGkHJy9nKfydfzLOhBhcC7OYZi6L8oezzxMToIc6kifth1XmzWs
3wWF7ulicOMOQXmOPFK3oZLnLE0GTJlOM8PqizIjoR1reQBY0fMdJqXADZO5Imzj9O+bz0IAKXPG
wxyZt74bBclNc1/9Re4eASrCDPI+6yeQU/rAXNod++iR2A+E0l9DrAyUOJ6oo+ooJ2fMQkcpPQ3g
dUswOueSfA1/WFUA2viCVzqwpzwh6QXK3egsKkaFJL8RbE0uh/qY+rdsOxeNVf48uL7N5bjhSiCn
oS0MrM6TxrbiwTLNAoImKtwBVql/mIc09sV24t0DfNZ0qBuF9yNKmuQ9qH5MemWzrr7WQZ4nNjXO
YiJYLDWe8kF3k8MUt+bh+ijGvhjN4nK5QdQq8EGCMzjhxDyJxK7ZCBTvA038lVH3t2sRT179/6HF
gdva5vgs0ZIQYI4ERJGj/sMCfO9StQ75arLnIEMFoceIM4BOGRoyt+Y2YZzAkL1QUhiFdQNOrqkr
fvVI9wh4kLdkKdTqS09TlCFgu9GtIoAfT7n+iL+Cj6VAv5FnP7d9hc48xMrbeBkU+578ayAp0tQa
EkGAS03PnnGCQs/lWIKM70N/NNv3ogHsg+9aqrCvKCnorSuHL1osbE3Bw3IlCz/xMrKfM0NeXyDP
SLFD2ZM7F01s5I5cL0P90xo4bUCX/IfDEKshbYfBT405CJ3qEXkoibwvJ8VTjk2E/eBUH+oIRRmS
MHRxhavoQactHV+Mb2GgXiSHpsln+TFqzmP+rD1jAtlJpd37KQDxmqeEN1JHbLBLIcWAaoV56FEN
HNLswFwk5UOFaM9JLWFtOHeo1XVXxbvXnb2Nw+ZfwiOP9hAwWDFUeyPwzFJmadFl0YVJrgHOkEen
pnSswhjHmUa+ovhRX8Yi/SmLX09jJnn4TNVTnZ85lFJJgfoJrIT/2uZgstl5CReBYvJsP7vqyCp4
GRaq1yz4tkaXqQsDLyMys9fg/GTGhKMdDOW5ZN1hebLbiu4zdyYnyCitlOEZLyke2vUjCcNsBqLc
+rz4dpx+UrKMwA6YM/ub6kPQKi60m4FipvfiCLJ/OKHO8miWfvFoVsnCMkpv7h6vyxyVGR9RCux/
YzGbaf36EbcK5uqC1MfoOi2bcrjSPWIBc5/b/bo1jMOHAToaE/Z9xtWeutRNgp/PoHMqiCJExQbX
RMD8EsZYDI6zGNFfNTTCwd3rT2V1XA/cOJbslPZBd9Libe3kjkzwv4b4NraoZmhwFh4XA++8iWjF
A7fFNw5KP/wvezXRhrCyuQykf54Uu939DTcZlE9zdL4LsFLnuGlZYMRxTDO9BJEDD63yBr4iKnPF
7/erySHOGR7XOV89fS71gDC2Lehxm/oMZ1Z8N6zpZtmqMK17YQFBXM2AI1SrrBSyazYWsU2lgYBg
ATyWUvRHRWWOsbg+YIRbPLWjrJ9Z+NRfkrmhmThWQESA5ZiuC/Q7Wztomf0YkkBJaZ4NBs1L+aQU
cE5lCxZ5cYNxFmoXpdA0yAVMernwWLu4VBsSutpX7ZJtjwNJ5JJ6BpoEY9z32MENpew0wXveBcoU
dMdYfA53BYjcWIV6tsk99s0p+BgQms2I2q/msNCNXok8R3KB7wh2fhRnC1KwcwWJbfBVtzOrGVR4
wY+9NYX6P4gCcQL4MjeKYlKzOSsbmcEzz+QSt7W0C9sBZbfWCdBm+IR2T5+J0AI439GEXczwpF1O
4i+3BnhIfIZOyQNAbMotzjcK60GHvcwpeaP3+YFIv9o7fhjKI2e3aNpnRSlMCdLvs3sigzJpMxPJ
s4U+QBbbWIIE4T8tXe4VMINNiibr/0ldEMw1zQFd8D5LL5NWk7Oq8TRcnxKbu+bGOnPb7yR3iKf4
pRpvdKQFlW7XO3iadtAbqRBXSl3NuBA876F8lHAXXZZkVBUPFZ5p3a5rN44CG9riMZYW/r3NRJHC
okX9o8gIZehmVmjwgYpBSIoU+jdbE50w1tSeO1TOgb4XfJzhJfFPd7ZECrhUCx7BdNjSTrxt+uHP
Vd4wY+GobJ8U0hlUQ6b9bT7GR/3M5GG+Otc8sR6oJIqipkMuLpN8DpqnewrqwaXV02Csh4BgXSB+
AoM6vxJIMez1LCdXnJMtzgt6+fO8Pj+6CKVrTiNACLlzfFRZHPgetrtk7K/q2bpdRZWtsZ1EVSbH
42S+ghNP5D0pDnrZ73QKldNuAOpATZ9ShaXgDfw6Tq9ZFNjPUNoWx3iEgmBKuHln8YPro4sOLHul
kjpApxbhe2i9Zj4uglOtcdN/1T8BOpER6Sf/m25m9VpQafm2lh223xzinpWvM/sBMpEidOwo3Nac
xejSvaGpcBNQcQY3S6C3tNASAg9f5Eq2urdzYmD1Bnx1mAiSlWm91kUuI3u5u1/wBlU6GS5/VUtV
3E7Us/cr6XHBDLYnIQEX3Dj0p3AuihUVAp0whOMjk4jgJ3dbPOuXQEA2t2THZjuj0cZQIVBEEKjy
QTp4RHnhXAGoubIQEhsx562w1xONylTOYEV2kVRvH5cZ5yxqQ62wN/dcxUTLSyDPm/0CGVK1DwU9
IVzt57eD6ql1J9hKsxjsC9gKUGxG0Pq44tR7p0p/3MnEKvu5Q/0n0Rh8ZYNMByODfwiawS+Y99DE
tLNm3CTNviAIgUAFCi7NS/7pM+7oh4UnKX5j500E7tYbWVRsqtl0jGjrR86Xdt+iK9jEnDox4ehI
Io/Dp7dONacQI7iaFTyd+rRQ3q9AOUd2RQB099a+LmOQ6GtgzSBk406G4dDO/RMJ2Ef3tr1clird
5dF/X4Pd3zgvoGwc03AGeFByv+Kbk77Mp9uuyasizf1/SofX+jMzW9tP3lhcbP5hlUb0cMY7vQig
tTM54UYC0rZ+jJ1U5PuIVH6WRvA8B/hjqgaMIFkn8vhV0hhvVz05UWKGhP9DpIInFnn2RJl/6XNK
tXAwvKRdRDlWa8WiYKN/cAjh6/5jP8ayyFBmLX64ceIKv0CIy2675PC2ITIDCTO1mQzOW6UJMkbz
Dtvw4qPhFCkjn5xg2FcIqvhRS7runwfDa7U2PHS4yCOFHcWgllGPf9wjOGfCxAUglQgGxvM2AT5X
6YqCl7m2fMLSU8nKArRFr11WNzfNV1cQ+NeEOIVpRBr5Cjqx+LXn0Fy5ZIoJK4mQaiiT7woExVpv
DKWYqEHRqsApbWXe02Ilumu7jPnTsoK5addDAi0hszpVh3NyoZWNb/cQmdiaKAwQSLswvZsGCbTP
hpJfixtFHNfLfFjj0mF2A8v+gMS3Yk4sMkgJNtyJDWdUyJTBddIWWZBIi9kG9MMKSi2atDj7cGke
o4uL8jxPDhgxIgvZ0KmdXxCizM/k2vLiRO7wXZxSkkPDYb/W/c42O+SzcFwOI/wkdKxwXNZkUnkZ
94+ZL52F704clK0zKeK7RgxChE0WJhtZeXatKtyPUxn/hi19rKbsuuKRGAqY/h0UwBZ2z/Y0NpzO
8RpXEDkFHnGwPHyI2tjlz+I9kNCwpI5eBYn6oR4QzCv8VptHKzKcC3gP0ZFpcTUfVcp/BgLX+paQ
JJVmNVWQVoVk/7lNEOAWIIGzztSUBWk4lY8LRHmlx31n2oQhiu1i3ugOr4i+1fsJdMkowM6zD3w7
apFAJ8at0YB7OLwQ1XGvrPxOqGxK/flFS8hGfE7xtsxE/taG5LXd4Fwpw2pr7odvyHHNmRUxSYnT
10FTy0JbJatiJC35EJtid5dCt0MBMkWX50q9150i/C7vJ7VfCEq3LIp18jmoN8ODH59C/RozFdlr
snq9pSxplRpaCmEIxtq8VEv+rFt3UcOdiVpYLx20IEWM3IXRJP87r5xu0GmrKzywO/4mbIoRcKHn
2cWQo3b2aYhy2F3l0lk1l0H4qQJBp0fwi9noxlYdPmAkmNtgokaOo6deQ+d7pC3iRtLDI5YttiQ4
xhYuuHZMpg0D0+IdvVobTKDAcg4G7mIfyp5++6kVxU4vHXGInHuNZxtqcd8e2+UWzgs1pHnDMPSu
vnbT24cSh7ppHjvV32SOLpZFG/QWwzOPPeHXmn4rLAJRShvA+sznZASb1OjQSOjLGmfQzzSYbGiF
JW4xw2kxHjIUCEMvk9mHj//3LBXztxrLZ7JkwZCDlpt30UX8LrJAjkHnlyyfQ9Eo5fPkEMOonjWL
j7FkN5g1E0/kAtypz84XCyOR8Vrs1Vq+GKvROukOLDIHATE6NCoYhns0+Has7/smV0Daq21HHd1i
8gzHpJjtKeZYTIEWwipdZHJPQUg+qWY7S1FjGdIebYLphKesEuG+fIHCR0sUL+2ynFRX/relC2v/
0M4YjnU5ca8JoN1ALy0o/pjRcKTFHPmwvMpkQIoSOjQA1pcTQr7ZvfSndwEeA2Qc91FwuS0cSTuB
5RfKjSCQjVJMAGObupeY5tQL6BSt/vOUsbmtkp07RH232/W/mpZF4ljAk7gqNjPCHPx7xuGDjB65
djysGp/NpvMXE2ihAx1952Eiik/Mrw1OYbR5f1OskVkV519xFcXgOHbFhIVI7c70P4gPhLauVTUI
Ijn+SgxexRw8thYQgo+LU4F0AkHOlpjgzeBrTPQbuE4BEHZtfrXm25uVl58noW9wvFKFfpdMwt+5
xOx6okS+2upplCVVGiwDn4Xgs2FFHmEoZvdxOaGP8xhBOdDiWr00Ai6EnQMERwLJAhtEGWYVULQ8
MTuyJbeYPZ9VE7tb7OgDGsnKsoXSiqJGlm0jTZDnp9gq9oeLu7nWivDIDYatYv4N27Cyt6/KOWri
soFbqXjGG+MNvyFrja7YHRpZTmPQBoY1ySA1roXmsmU6OWqnBUpNZMQ10cnmGy6ClR6889Cdkxg7
Chv3ifL7Y8wqPEh1HTkUldUnhqo0Vx8j8LXHvrOYYUUtPFp04ITX4HkibWiOlGUvWTeLa8yPCXV7
MytLovVjPQcoXYuZS2YSijXmlG5HiuE8N201IoljppIwJIOzbbrf8uRt8UywFBPED94KJ7y4i7xe
waJsHqPglPqzDn3GA31QDXAMWk8EX06S2XW7JeaYFsy9wHip8qPXoKmqcllBFqHSEp2R8b6fMXA3
NzLLqVvkIiFnaaNoCfe2t35crEH7j0xTjnBKWCCU6zaWTLYVUFbGkwTlJIa+biaXIO+3jazbJ0/I
ukYAH2OC5h3ljKnpoGCl0EwzxevSXwqFeA152ZhUcsuD6EpG0bBN4oQ9DseH+AfnyZz9Qx8OZ4Lh
qTC+TT2S9klrj8Lav4/dIbi79sT/o1kdC9+3i3VGisx8vJxmYK6hO+Lol6JyGr44FBbP1BjDdjSt
Y9P1gkhh9XqSOIzm3BAEDMbL0h0jHc52eB9PYt+suhr2egWTaaWjF+aHBFhIjq10sCyqRW+LTj6k
H2Gn4rPiu35xCbENAG5Pcb0GjPumZ0uuq97abtyQOuR9DjqdYLkd6IFMeBG6SAj1fEtflpwNCo6W
mAw0UIWJdBaPwDOSKpA87aD1psqMDemqmHC1sFany2PxQ3KmYr6YPYXFm9tZMqybcW8766eq9GDy
Nmz0BTRlPO3+Fd3b5PIyj8ZM+b0D82sh8E8WYePWDWu2oQc46zUFV/gVt/3BvMZYYqi2CZQXef1R
f1yVthB8+nnEnUa1bC4LJoxsB9TEtCYM9kYnFjRaRSK8P+kxq3/7/un2xQYmABJlxaLB1Htg/w9e
S3kslxnw5FRQJiYotIiTBGbfjhk4iVfvwdVc9kRIAVxMdXSrQn751gxAP0OPZAnpuZYGdIjR/+7q
TM+dh/vCEWCTj5UfV1ocJckkQIt2S686xZl2xmjamsPeHflgccALpMoi2yoj6EoYE+KQ8EtFT386
DC8wGJSEHMDzHJcPlQlPzp9E5idhpyvt+31n54gJ8Sao3aYdGmV1uc4Ov71OsBq6vtMnttRAg8p5
VLopReo0Jmjh/fqpFECj8bB3L47+wR1DqXeNeHEQPZyi9nF6zFAgIJt5wHjjoGl+wGdq3PbYzdOs
KrjM65w9iNU+lkCYx7HqbyCFqrmE+R/UEy5RggMI/PLvG2EkGqqHDm27DbaLlGezhf47hm3/2YkW
qOQsutyzGPRnxQFVCMnrIJd4asZ3yd/V07Y1qvc9KgsQv6HVJgb4IttidR9grBVhB9pLep6z9ym3
96DAt+m/R4r0d1g7sOitBGZFx/ZSc6fGjybERgNbyEwsnFlFnrcl3Oeab3OuwpK0flHrEXAdLfBV
mVoLp29+kGCzlAI+L1hu9mAMhXoR8XxntVsM2q+aF1X9nWiZ2OOSekc/nia+q5R7FpscP1RZ+hDh
LqDmgapz8t1c/JVZKNOka5wDvtNQvx/EKos2xdSQKV5fA1nJrsIl2toCNkeMXy6/VRtDZfHFqtGt
7pNBDB6mQUcpYem/1zCHrY/ZVmoTWdP/KNUa3DwCCZILPxdhhLnnU3Awj7GIBfJvYdRovJ+PLehi
bY2o6Q+Y9qSdoBvabvOhPzaEJ+qgtJ0VTSp1D8pUJrRDTc+7KW3oSAZ8r6Wyl+OW+iHp0Y/km4ZU
iRbPPhH5Na+6G+00hffJ1WTovN7PqCPmhFwSARrmkiXzwYnrebgATfgEVaCS5E+KZ43GT/k3LwQx
boemoERK7wlnTfDTwcI+y4es2aoyP51RsxIkKkXC+jlLFyRPl5L/r8tV6ehmT7LctyBRuAPp6ZEI
LdP/a2/JWlQHTyy72EcVeIB942ILLtZYgCHi8RqL98pp006tohuCNrwAl78uyxMKyjiUYXLibyWU
p+O9Z3tJNN4dJoh8CIVus7CsaIK63u4nHlPHSPXQactAiIOOWhaZ0rpxaCVYb33jgm6YDjHoFOiH
dl2PQK1HrEtov4e5ZYEHORPDb0GbKBPPPChOEe8AqCuQ8BXH9HhCUtmKQ89unrBavO1orSv//AbP
ht2ASlN3Rp1YwPcfM5Jxlr+i73MaPHiXs5BqckpcZw6qpMl1kbBKShrTs7xSeqZIQns6I9FsSIzR
1X8TzdxZbtB9dQxa221ip/P/CG/YpFRxozON0Qwdi8KVWUUgvzFFUWyMfQXGGPmywvDgIgAKCGNC
AvbuHbuCBm2+6T0bGtxvqZVfeuD8hBPLkNsmNW21zQ61x3aJy7k6fgRbbMTxXF71QQx65WqqB1QG
wklHbifE84fICHTqZq6RF40LpAxHPyNKzPd+AV10yHS7OVwcHNT0/lWTDUJwDVAj18tBQoZntmxZ
96k5BWiEpqdiIH/Jnn0umsx13IVAP7WhZm9N21yNZ7r35zeQjTYCZeo2AI26iZayyPhYNpi6VBr6
7IROH3SenxWW4b14+7KAu78HSYBU7d1aqpvGjjoHLS8qoXyIPHc8fqTKGZpF4XQcoa3wSKV1hJTF
CC5WoGC47C2tIEaixssd79HnEGE4o/kv9ioF42HdHDOhxOAngXxNEA/AaGBMCmNcVFXSQwXw4A3V
eNq2npmZLNyIMeh4xKLWeK/ZILMFH8Aa/98TnqD64CHQlGBRcNKX73No9dpAwlMb6YQA9DyduVDP
FmDOgFezf6s3C/QAWJ+7I6fth3r8ykTMo37YFrpI7Dt0c6mj7lIexzxyUppjVugusiVsQnby9lqv
IF/0OXYBcq3Qexq1VIzVmOs1nWtdIt++TylDpvIAlArahS26wxNkSBUr9uwSoksVGThYPvttxDPF
cPfDs40cT/pjjSqJDfvac94oZAjXSF9/QMq/fQEVymBxUQyY+IbHSC52WOr2eFa6ug7JYZjy/DVD
iZRATlFo/5w77UPhajllndiXo0RWZ2Bk2aRALrZqQTecFhEHmyiIGRP8zynqc+iNZVrvJFlEYBv1
OmgOswTzN65eQBt72CvCMnmE4HxZpYAQ7TUplcaBSIJ0wW22NI+S4VcES1X9CbtMPER2PAzhSORE
Q4K/BE0NTPatrIe1RIGsMWqW2Lx3VhZ+cWScB77ZNIaMj8q2hXZ/6AFQv0MQL88mfM2H7D0f36N8
yJYIILqkResmJM10b8T8uDJDV3V6VJRnBK+3glx0QabSHDGQl0uN2TBS48aNAnNqWr+K7XHK6YS6
9rUDbadaa+iq+iq24Q79/3QbMikDVMY/rVasTSTNUsVszNxMM/5Q0oLwbVSDWNN1H12qcJJnCjSl
j/ZU/vgtxBMcl3Npi7GdqJJDw0zNu/yWaJl4wTFNFDn3joikZdhJWNskE1H2g4caXDHWeRrqaWfb
bU/B+ArJVBLsvQJbhJWDOXWTilVgvomkcsRE+wolPRqlJ90QTxmIdWoEWkbB73OPey0D0KRSR6rn
/PyFPcY4M2movGxs6DEVXQdZ6HNcoka5FookgjH54qPYh2rrlWupBmTOCxvCFd1agHn7ipYKTUOp
YptBU+92KexW8jO5jywfnPBdLDiqa2CphWHw05h7HJRH8OJfk4r/7c9m13hm4LhNI6TPcrnbqeId
obhaqwI9AxoSsdRAXlal8tUHMcIiP1xnmq6oC2d0npu4j9MnxG7TQKn2Dt5dPz6GukToyM3d5rnv
Y62cqvSurs49zsDb+mUuJ2m7nZ8drS3nFw87a6+Wenxzxf+HLRRhBySY0lbkf3mqNcErN2V4zTdI
WIUp//kvboa4hMZGTYgc+puRcB1gXouSW2KePvP0vJLwDDn3k6CW612v3GhK6LBwmfUhjr40IUu1
RBprZErrT54AvoovbaJ+D0qnUdOAaUXDiz9fprT0YSu7GKXoYEGphymhwHURq+47rDtrKCUlIN/3
GD8WiPicI8dki+zazL9bKxuQpxl1BVoZy23wacwWZwQXMyM55bGLqwHvKqWRE2nEAy5F7rFoEm/q
xexGEwSuJiWaZffahcwO3z0xsjL41maRuoQDxf0gb4mEyb0ZbdnKKmuSMfZw/EHi8VLM2P9HkmIm
k4WnlUWzGF9cWyOysuwLi96aiuTpRzOIu88zydryh/0+YDwgaZ+DUbCWf7LtS/PtnYp3x9O1IfW7
zaKTnyfJAyJW/Rgw+ptQMBihqMTmbWpg0cTlp3h/Ir11Hz4aTdh/qHypV/j79QH3xmkzCHFeDA9n
L3veniQiNvOjIyi0atmJ0WrGTNepr+VJmKns3GXPg4XXsjYTkZpwnFCiBq10QMc8mbfCkJmZutJs
XwDweq99KHSHniLsjFedZ1qo/xMm9it3GMnC8ArBGHUeblRaamFNXe4riFel8wN89115+We0Ysvh
DuoDUpWzhI+2E0c2Z7cWYuUNd8+B1PrgrW09xhSHKaARe/1DWQGu3IphSw/o+omvieHmFR7JYWUS
/Bjp7dXwiWTCn2xkjWgb24wtMNB3WkhOz4jPQ236ww+MDWrAcXPbRaKgePDPc9LBg/yLMh6Du1O2
GVijbHyxxpYBChzA0oJRbj62xkEqD+8fzEbAXy54OAW4n5gcytZ7aa+x8X3X5oJms+FEAMyIDXsU
tC5V35VvOJPJdb+p73mUTVVUtV1NX52r5077+qZegi/iU6plqA+FZU4UHPGqMNAka+nT7lDB5Iot
nVr1+m23CkUTGL9wn7WR6S/Zq23xWJmQi9/BrTdoBK9Cq2QsXDHuwQG3WkrXERrWya1epO8jZTgm
HOMuOn1VD++9qtaAUc49SizEJsT4dI5CdvSVfOGCEahsVRg2LMTEjDiaECsi7CEcoIPrkpeSDLDq
ZwIzs2ZjEEJ+PVDtshM/ieYD+aVOvlPHPZcWCQeWVEoaTRYIe5RGoQXoZ820JO7E3ThoLJ4K9vFO
YEkgFpajWuak6DjLgcEEAezFAxy40KzV0qbGvR4OvilCKOEjWh0+1XuCguKU/Gft3lXbE7Nv8vvB
Gf2Z+D/y9734l+nTiMQRj9O3cvic+F6U57/J+VeScVSDcQP30JgBo9Vfl7lsKIL9G6GnD01HDAFx
WpEDui2vbqVs8F8KY89M+T8BgSKlJoRJ2Tkgqkouqw3QYlMjgVLQStpTc/68l8lFLFdw91IcaMrg
Sv59I6OasUuS/AbaYMLEj64OZWyuOJirPNtjhlxxM7Ua6++odO7toYolnG9qtSuVzPydWD9BIzTM
lGh6oNCmkMSL3pyaLAUbpVDm8v7WBP+IsTF/89R6Qh16Wq+4i33+OgCqTDynPhTxZHJLOFwh/BQt
CCSaK4efB1AzDZMuKOL9+YA8SPtdDRzPLQ2oIckUqp7Hz9PpgvUf/DG9QpWcf7E3ONrRztJeDE5l
2Uf2j2LdcoKcVFCWuHQ0TtE4NML5ucCH9YwBtOVvnHQI7tSMLsDdchzhWYcVBtlVsDqHIhwB4XCa
FSbBj5kILE41qkKoptUqIBbvd3i5KKNDw/78fTYT/P7dIcTRheCSpwsgqsBChLEkvxHxaKnNBMbL
FmfouOXr3H51L5uats19U8Oq2cqkYLI7OeziFZBF/KiB9PBWMhH3ynoAqF5zXnnp/fg7fbkH+/L0
bN44ykrcC7QJRIsO4tRvSLMq2LfI8PhCVMjuKHzUiDEB4aH6/xjA4f35WeU2aTMUdosYmRCcGBVk
8bYq666peAJxdh45RFsflbY847JD0c6GPJIbrOIAPj7+nLMQXpIkQaAJfEg6dQXFiyKgeTYMgdfD
hO4X0+YD0WKBFls/zONoLlvqyEupcTrMscadEJ57JG7nNh64LYG0f25EvEwAoq7CuHVm7l0t1CRb
TESdQ57p2dG4UcXjHyuMcKPJWEmIbtlJuPQIOpgPr+xqDp0yRYEMBcT6J/3ABoVI0Hj14YhnwpQu
S6rh7E+sk+v3RsF4i9h2Uylcbzn+kBf0tOOMEuCzH6n4eWqkgLHijTmC/daKLbZH31vJ0voS6YBY
mfKhIXDBfpXdzY7Tr4xDNlHOfgq7Qa0mF7y76S+w0LrUyF45czPvJMkGOloDGh4DdQUVXJYHch4s
JBFxn9AH61LRAH9c7rCiedgQGFkUfrRjCO5W42j+GZYm0HSWU0WrdQHOSc5TG03D31+FnHtI6zEM
fIhmPbns51DgX2ctsvi3UXpS1uFfFxeaz1+EQq5nj1rP1e7PcsgqM6APaEg/b5MDbmpv4Hr4teXs
d/3R16iTRsNGfJOQFgi1q9OebtvbG0c2Hi7qDGh40QVYwKhiz+62x33Pkww+bTNmDN4thxOv6dKn
YYjTU36BwQh+dMZGZYlVFXwv6VZB29GofhRZIGD3fNMZbgOgS2w7rt+q5yYaFFLdll6qERRsRwrk
hOpunR+80jyp9DuqsrASnhEksjTD2deoUbbHI3LBcUrL9HwxA8nU8XZc0SxfZEth4A3la8wc5s65
3XCbvFiwgMR1n2ss6Ft4bY44100d36XuvPawrazPrwZieAexpqX3vjpowLyTd2oDHijIwCxgJ2BO
JF6eHfob004enH83ERrjDdlQxaIy8bXICZ6LeweOVSrJzAIe9k71nlcosytEZZPepb+eWQcUlFVJ
r1XXVCbbje9VNbxGQZlHSEG29aY7ieWtvNzzjzgmHD/nx+2teUw3TFzuyGsIWwYNWuEc871men+5
L+dM7ZvESZnMGAlYI/gAF9CIMUcZTdpncfcmPYxQsFdduTXl2fSKlm1tp/YiCxY6V1y9/FU8iECq
Pro2j2bXIr5JjSyFh1L40g6a8MAPGESrc/IU5OU45PP6UQzbeSn+agUsb0df5oyTFnu499tHEuce
QFspZpgGPM34o/pB+9L+7a88UPJNShxWL7ZZV2a3/LEtvH1tsa7QQTlzE+BdVsZ7nAZ1C0HqKVSW
g1crvpAJKcTONykLpCeNBfuLcalF36Z/BMKMPgnGC1NgmKxwcA4rDeATEfZswMikv9M6tSf9pCSY
g1BK3JmprRna+tKB54S+07pKnxcuOCDHQIplwNvhs3Rr3O0q5JsFKKmLKEimGNQkbPY7gC+1Vw9Y
+eX0DRRH+o6OcA2X5EnEdGf63EbJUJCz6IKQSo4px/U/7hET4IbcLXjtRY9C+LePTvNni77bUaLj
22ezoqAvpq+W9pfZdAsCr/WxTWdP78sYX+Wug+N/+L8OzoG3aZ24lEShSn7B48EMPRTSG60I9Ptc
v2R8E+J63NAbdw1RK2BWXFJbLvHE1nOF2ubWOae9uRhPCA1GvNCR0TafstJ2K5e0e5i9LPtrvZsd
y40sbABF6cqSveFpaAWnipMAz5pfZ73Urviafx1WRFkzdj2TkD2CL809zY6eR6zrt856Ll3HRI13
EXNdakDTIJ0raT8fzL+ZCRabtp9PLN3p7bRwAMLVicI/VwqwdX5ykzj0YiipdqcDRy0X6iDOcRgr
5kzdHxHJwjGy6HiRlDnmxNTzT/BC0RW0XEohRQvHboxyyGNQ5f817ft+d88ti5WC7p7CsUoQ8V+Z
CLT+nGslglbS/6sB/lsrDlG77tYNNinUKQgnMxRfC3VUS4mO2qDpsZkKDODwq2FOTiXGNxqryHlL
ueMsfs4eZah7Sv6r7iZliIUemWrz44szjMlAQjPFtnT5LLai+E/vx2uq/SB1W4Zvnn4FkVKU74EV
EM4s/4r2HlLw8myAOYQWtYLSUsoRLuZocoaYib0UXc9mTvzP2Od2AvaaC5jEC82B8ZcwnGhXsw/8
OcKHMvkQq1kqLKgQNEs81WR0t7NWzrVIjPj2VBDyYlfkhPUwnTKLciRi+yFEg0wQnyd5QvIhPXRT
yclWjQl0BRj2g8keWwtNK0XT15UnmFG3j8EaW0hV7HN1+oXBW81X73x5PsW26ChpINptYzd74Whb
ZJjb0eEXdhM8UWeXJMW3+aqINQ+2pyR8iL4W2DB1zvJl34Ds7A21iQtET7JyaP9TaXBfpWJOfTgL
2x6ibTC5B5z7izkjG1cVfolKXLCJRDX4JkKm5YWr2EVNkX6nK8Zk/GnpWEON+4P9GJAa+7DMsDrC
zgW5hM6ue/bP9+IrhAWF8mhr2LosVJ/ONPFLgOoRYpZMleA/TGkmqy2JUUCATIi4pxdFwLAFWusv
wLA02JVKFgHKgTfaalz0Nsfy1jHqQiH+bgwbsJJTvgO7x4+1dTQDouZ1Ydk1SlGbaye0zzW/ybFV
BhRssdiJFXResNNSeCmvNBpuYRnaOnRN1I/6twDALCOfpEhb6tVuJd5mVYpnRBTr0Ur1uzVn9l1X
MUUWHOGbNptT0ch3HIro/HOZ0DJhH4aDGMqjpdqnxF9VpS9wCDg/6B7moVpl7DW80KtyI86SOKEK
GN5+qjAULZ/TUpxKpmUokWm8vFu6nG9tERBZzhA+JCdmpHqljMdk4NbixcDgJbM4IMoecXp1FKCb
xeMqV9SPTPtTdhh8O2cKBtU4BdzZk5avv3rXkqtTULQHw0r9MZsW6v0qjnU5V+XEJ8L2gRtp3y/8
HJvE3fHVsksKP0FoT4qz0FVhpOKG2MsmFWA1TG7jXoTRawDp8jTOCwQunYDGAFySYg3WmrI0osPT
iYtuok2PqGBItrSwv4UT3n+0BItaVbtfB8tOFUq18FmhRAQM1xc2j/Z/EwsxZyc4qsX2WujX7HYJ
sNeu5psLvjesBqh9KuiQDgmvTXJqZwa/xGcKBfxFZ6kDDHV0XlOWXTZTkQp4SybwyDmH1FeYmC0j
TVIQMdqdht8XsnM28JgIvEV2SvD9lVCOnJuHcZxCFVKitG1vZ5NkPoBAjTpqdc/Ofoomx4Rlc+6O
QDSB6Te/2K/ln4cKB/8KWWVLvJIzO5WGSsyni9spQWWHJ4pIV5Sz0IcodPZ6TJyZOzDAETuZvx7E
yvckvikB3W0X42/qGhMVSalw7UN36sJIGsabP/a1+qqPx+OEsOrQnTg+UayOS558BFZ0ovwkaKze
xP50h61rxcYRqiUlDUqbwUCdJjLfniEe0X6Qg5ZJYvt5tRo0Q16fR++8maF9PxDgr1F/5IGW7Rv9
Z3PzAE9u2gtRNpm/iPjpEW7LRHm5Yiz9J83BWmAR5m9iPFs/veM/80uos1UDzHzY0cXDbB5j9PbD
6FovbDclI+wF6QVDWh3hyegF/oxAuEWEmq0KIRTOiDGDEu0uTsJiGZkWtoib87mQ48ggNB268Aij
9hvXEYMxgDj2dU2Ifu3E1WNzYTIimG+SPqerJAvrRG7Pj7dMT+V8h/qB3m48lIgcZAa5zfThw3OI
RafyFpQuuy6I7h1SluARF18yxSlxqHh5GKjffcuvHS1dxiJns6ITYNnLcWPflQbzTgkwk8K78Jxs
JtvO4+IjHdrrgWwgU7StwDtHiHniel7G8gf4aJrKdXjbnr9mRq/NmDEvMlwsyIuZ2R4bmnD792ra
icDUUR3Lkn+lo90Ie2pdlPw73ev1dJchQ8APvyy5HnCsblQlxrlsSCOP3istKCRrsNgKgoJONw9Q
wjf5/f9EI1mBgyouUyFDtQQBG2QSgT+YF4T7gEcSqnly7MRSMcvuLCetkAY6+Go/aiFcbp3zRYIx
LXYWUsFaMCZop/x1yivValFll0TYdQ9RHb2q8D2LuY92DkfLublFC0U5OeePLg4aQnjPN1GT8Oi7
5nQY7G/SLg6fm60rCKhGWF7DPLwHPr9blFv2+Tr6RW6/bO5LEm9ryDGTnkRsRI3Itc2JnscxkxCV
kVjc7yH9ErmDjaip02KuCdQBtqdK8ayAG7STPtXpTIvUbtk68X04BzLcNMIeW9YzmFUMaU8z714Z
WKVzA4CzDeSdBqNy8LvlZJv+f6DdqC7MnexuYJkpclJEKXVp9i/TiRPHq6i+8k9m3HWcODZAlqCg
LVn9PPsRWmce9rrvfIvvyZWUr2zEfq3xkcDnyKT2G1C98DkWaEKkbap3ztPnYzjvojHuigvXpZ5q
WWPZ3LUiq+L0EYhUNIQdYSmjqsGbTfLC4VmvbnFiwjcMPmExg6vQSWQz5kHy2eYc/1+dER2Xw5tW
viKiPFHOIY5ZaiG+LnGzQ1ZkJZIfzg1ZJmySne8ZLBIZvCLr1teUDvf9WvELFd/pwGmFQhtc0Far
6APtriZEJnqGWgzM7ss8Dt2S7eKVRqsP8Fq5vz6TlfQ82YJFC8Fq3Exg3swdbT8OQkNx4bETAFvm
t8MTabCzDFhE2ddBu2tEyBe6bq6aRpHyQWi8ZsO8Swpho2DB9Y+SQdt4jphgYhwMxXZCA2TUYGXf
DQJ8+OlauFicvfFLFY2fIiE/QOlnKw2e1xSvSFGkK3Ur6z0JiuE0e34YbamHNJleX/RDn73nqL92
ulI5xk/BKsPKIdVPNdIUqW++m1is8eK5wpySPhNKlvl+wEiHmV82QvEOUSycEWjMXB9LGN118mhd
ALAipDaLpFYGt0hBhBfLUynfJ3bTyRMr6hdXdgKxeJRmwJ0RXFK9+lB2Lm1GD5QDTpLnyO7w2Z7d
VbV5Jzjc5PIn37P4VebMkCwtkMlHdt2wUBammHz13AH1lEyTR8GXrehPssR1eGBmSwBH/yZO13Wb
NgZ2EucepJmKoBul36sWXvW7RFt4JqcsXpvjH2YepLhsbUB8jcL0AtrRNXbuokp7VINRhhdKzHjV
R7VLDKHB1Y8yn2uTns7ZL0jXu6lUvH+rSWIU0GHN8sEZ57xZp4VOJrY9TGoIuUoKZg352VVObKLC
BGRjO6Bk5EYsy93RUh3coDpMPEM+KvCMsx5eF/lpsOAL5qDLegGQeGwYJmay7bcE17/vppUAOY8e
20spLQxlJUDvk1SgSvikzQ9PR30OpcxQ9jZash59x19keOX4C9RzXXCV1yzBUdmNGYZ/G7cI9iPM
24k7OJl/zsyn4v3ChSiBVlPuevrTHxbAcUkXW217iDXLPsLhVeHsa2Hcgk+tT5rGp7NUL85ihXZt
4hLfPtLq1x4sLv+vbK/IILUTLB8oo/bTmwOkTcuWKLH+gm3rGSZp08gbKK8YUhZ8227d+PupH+x6
eqxV3ZfzwhnnzIzoiAOlXR++ReOAZQlOeQFEoH62Yl/Tme76rLDNkUyh/V5Y/z1LD+gb5eBYB1O9
BoKrkfmU+6E4ZtWLoOKciIue8YTmnY1cFRkhW8xARd6Fh/7OMpBUTYPFZCjWHgM/DLelcAR/dubq
7UJYWqkO71XrXzV5cOpS+83Ew9ORkpfjvdE0tdrNPddBiS2k/vLn/5Rc1RtvHJ4ru67fgGIyPfNd
XcaaterqiEji90mpPs+Dw/jrBhzmwgIVEAeJMVLsbM+6IJlrIikzAOGN0qg392uCzWOVZbSN267C
yOjLHk6THS5O9JGwrTkBIUR8oLc71ide10hMJ0dZOxxiVFBRRT0j6sqnbC4tSKEbQ+rAJTb6o8CC
pLvhX2x2UFGqMniqWx2X+zZLVOrtd/DIOOBzEnkc3tv3mcnyu9O6UBtUfFA62u5R0KvfPR55lGlD
BwNJrcGrVctNojmatvzDIcDUbKVoAyYCpzCksV0E6I8ZxX2KC9pq/emlsfUgp9fdPlGqzwGYc6K1
lllVb5UNuYoXCp/cRFdavkwVZlH6BGJUNcMi0RrquSOEygDOK+utAU60fupc5qC8gB/vbqLEtk4e
LvrTViowWCBmPckNTRfuompV1qYa5AMYymkVhD8DojTXcwQMFlDkyB4RX2FLMU1XoM1LG7Lfm5dK
2UHW4axE9WcN72oyQ6oHn+6wIvN+hm6Hsf60Z9p8haBr8fYMPE0I4gVOIzNPZ9VaS+qFQFqU+cS9
M9/3RkemdfnETOFeG6aT/kwWXmJy1GSjDeGqydaPbSx4JYkaE7jnNsIG42nu9dIvVUcsnCCusKCg
kKKvudLtrLSoAa7syvopowFqe5vHKtR385EXKnO5fEIdPUpaEk0/GA/bDNJCsRot/78rxQwj4inR
WQUmi+IjGbuBYjV8eiBrwksuW/uLSLnmr8r8/UoiZaTwqa0yLuh8RvgjXFQ375UZJs2sedeEJypN
DhfSZFrOxVv+fqWCsyrCMhhdxxFIXrpKNDMyeCiHRP5b0xj/olDqaB4jw9uTpQsrOR3wX00GG60Z
wURpfzljoKcvdbQiq3Z98fRdU8B9eyYluKjhXwpletKHXy47hRjnj4UtOgwZaN0dmeJLZ3Gijt/e
da1SdphGY1EGHspwe4tToqxjzZF0//NVmZPNEd1cV7UXGn2dX1kzZx1VgnLiplANZ+xfVdgt/92u
zIthHRyUzHzF+p30vsmo3mYMiqy7OZI2dTrfcymvgyuc7GcbQfs2wgbK+CgtWpXnjtXSD6yks+Gi
zEX6UL3ZroAGUhhER1Wigi/USXU15SD2fglu4Feq8JvtYZhgyIXixHI0X9xXmBxnVmRCoywcMPh4
BNStihMyznfFs2wnPKb92mVgCweRZNJB/BzoT+TeI+R7xDYLyGah+c9+Tmcr8svrJ4hgr5PGZ2f4
+aPGeq41W8uzeXJO9o43clOwi4iLfYiipot8/S+fcGb1TaV7idheQ3u6ao3MvCEYCrBdICzwlDaJ
lHGI7x1sM/Ek/mIAtPfsZcLTDn1q6VLpWyhwVKiL3+9abCKuNfWJBKiDhaeG4GYpTIEKO8zmDzEc
9YqQTwmjbHtcfPuLvC215jWFvSa91uCWO5d9jSLk/TyqOq+43rKMTsA7Tb57q9jnu0E4+cLXQ19X
Fx/WWYPkziCT+0aJzvtxU+9pucT1IDmE5RGo96Ly6Mazv0L8ntYDsddbCemYXs2FJVdmS9HUmm9S
axfjbTq5RajwgA1KWXb0BzB3bPNaBD3f9G99dqtuvxJ4fd1f1kMr9I/ePalk7vUjAo52W5F54EYx
jvVSH9/IBSO5JkyHxAo/hw8ecVXfh9LMTBKLOV2rNDDOtCGZ2WLUB6k783e1nMWa1O85fdwqPzVL
xAR07cJkkqopK6Xxpj7/Lwyup0ewd6WBSrNifQltyzQXAbmUZRj1u4xliwWzzHlHc4kYolE4UIug
2EO0rgXEPvuSc2IxwajVszxyLhD967pYg9gzFUz9DNF3VzLZ18RXmHR6HUqrAFPEvgXWxb8/aGol
i+ddf1FP8DHdeVIsDk1DcGPlUngRf2cLFueDLGBg3XmWWGUHt4y6il63H/8cZ4TYtvnYt4H5hU1N
ctYZQ6Eu0+kJQvuiWd3CYGo/wEw451GjCcRxo7Q6eoSxDVRKL7ljsUSIH2rfAxpsI2uRMLL/O7aV
LOFo9BYJPbONv18VLBRSlbs7r4DGTr8au3ui0ZO9aWJ/zjok3OkJRHz6dTyIZJO77VabCSHnWc1a
jR/J0Y+vznUkTnCcFEu/dt0NymmL59epIObQtupQGRgYaX8RV6l23QukShxyg54guSdus6RhlGNh
1hpXDqqwSlIeLOb8+xpF4uGXWH0vzs5I0hNHy/9FtNbtz2en7owbw5UaxHdhGnTvRCB0/8GnpvYO
JYjd6aJyBcIkA3WeKwgnfPkoIv0sgtyQJqptlwgq7I3PH9JwOhhr3q8lERG5HOLPspIjlRm0+AJc
Ds0IVKRGvaIVYQh1eeIx4PtAWvaRb9ye7LBMv8xZlSNRzKEss6RTOU+2RJwIUxUYB+SBakg1ysiy
233rVfaUHy0utYcZJmcSOppu2piJOKYmzFs1XPV8c7D9gl1Qvw4w6GzncTkSExw5IiQoJ82SDoUJ
ffdIgSzi+jH637HgwH6wzthkhNgCkh4Yw+bUWk8udeMOG/3ichGyzDRxm+vixJqGNkZgDOWub9eQ
ZPAyy3j2Tpsnqova+jonbO4K7JslIfDilbc/IpQqHUMhHlB9h+kgPU2ejVP6tuA496EwFK9eigpR
8wRYBbRBGPctrPN+R4e8RBDmq8CKGY73iKit966EB74WqJA9ZAyn8k4GIdwtyMtrO0ClhGJKqJuC
inFJNexkOzxUoYxvMo3QxNoni15UMJW1oIwI88Ahh0VLSS+0mAAM+pqMYqKru4WmXniVme5d2TJq
WQ0WuLto2m83sDDnaNn5gcCVygg67lNigx3mTbJ40NvcnGwH6VdJzTynYxKmYjs8WCMI3ob6qPF+
OWpA3D1BJsmf4xcNbdDTukNjlaP4CzIRa4Nw8fRtlDxKJrcaY2HFetbN7i0DokRUsmgZ8ue08klI
ajXkdr3A68M24nrHS/Q7eIWuJAd1nwFXU7FPPXFDYT3XPtL7CFe3heBHR2/25+yCpV4OvzfJ7TWb
vmfasQgKSm0L/i2SJmCd6LXe6HduNYvT4TvLASLEz/8kye95K23q1ce6s0dd1cTn1bJaWY+j6wLO
7/7gGaJ6i1egZrL9kK5AOXNPhBZxE3rwrqHLTc8hJKjxMdYGy5goI9la5t5U7N7s/b0u/OlHOa7I
9Z7QRLt57V2iNy2iymzdvKs4uD9lqP3AtLtq8wXQKbERLZewJbBD3m7u1kW2l+WkZqzNF1PqM3PE
RQlCcUalecprvAcJDXG2r33W33D54SfHWKzSqep5p9MP7dkd0WPrkp6kIHunJ0QhVYQiIxp5X0O8
Km6JsR+zIeKvWKIMI1C67bqNkYTaPnfNm85jXUCNMmH/8U6GCD9wz7sRhe02ZaEzdJk/BFbU/0fw
vC9L9nuFQeQlmlY0ZxjZMVNd84OQS73miqmD1hjCOYfc78pAkbJ3vtFARMdseQ+MKDwtV/1Azeye
EVlUgOHJR65rQa34qK5KBYSgJ/xkq1u+7y4nJZw7NoktmdjUe1Ro4xhfXJivaqPuIP+y0EAnGAK4
dz+FmIzulD+r1633G1huRb3JZTIcmTJ8FMqqF35soARtZmSAHX5Gj+SP/IaGstOAoLY9AP7P/8Zi
OHNam02MT298ghZXOrzswaNg1qPOozb3Iy66XskprbCj/DIfqNtjRdgMX6YabDDMk67vicbynTMZ
WzAAU4wyREeZO3uV0iepnhzavNA9Lta0VGrcJ8RiOdjzmaa4IytiF2vkIi//EqPfIWh17AoVLrVc
547Q7Ro+G8qJf4qWreV8HL8BE5Znspvjf42gZHma4bfKYn/ctjNbz2T9/KN9Z4j4TLqJWTxCndNk
8Ab0VUlFx4BEOVQ2qkLIWAw5kj0R/WZrChsqN4fEpeL1KzLoWcXfqNanMFbcpn+hZpoOVSAWcYx4
mIUkrvQ6JmqWqad37hYXcpQFjgtQNIpdzoLfFTU3CJz671PRnEme+CSkYBhT1P0i+MQ8xwYPXDNJ
gt88GVcCTmIpNyQ/muIDzmup//iK3I1X+oB4Z+4H8ASqtiaabfWHoiu8RjuAUxocmgdB5/mzgB7y
HaxjTMRxrj1ovM3VAxOy1ZZ6EYyeFnPQA6HlBS/EUpXdCJoCXPCPWAfZTI47AEes3jQG+6Kfl+QY
Sar1NGr+SaMfxDIK1Q0MBkjJ8zoTZg2PCVVzq04eAmjkXpujEqPvRZkDx4PY8IWhCTuk7vGKQv+v
DeT1qwtjkzctg9N/gMA1tprrTXxUX3QsGDU0uFpY4h5tHEZIdZLec18pYvLGkucCu2XwIyUxyAec
R7XaQdA7U9r+IY11NBZ++tCjmPMY4wPqt+cA0zopEggMhj0KavtsKD3N4gjdPQy+lyKjEl6I99NX
nlEFwgEsuroeLF07uS7VSzey4/XWvcSMYD9lJBtGtrJ4qQ33zJJUsDKiSu+qnY6kE1Nr/ZctFX0P
T/ekF7PnVTh6z3wXlkKCvKOxyhLxikgtHnKOgAFgXkdDRZGj2E1jgM0SO7lKaPAXT1NMI9hEWppL
UQgUClMwubHbBxLZxVssLc0HD525VdOj736UHrA6rWH0j12zb6QU6nS61+uM6avhgOgQIxBrWL/q
3cP9XGHlINEBK4sCekZIxRdXfTqS4YPN37W3GgUFdntci0gdWLAu5zZnUwgSG+/B8Irea2pDj1n4
/g8v4zwg4rKjjnK9A/5Y4jjXsp7EonvQIp8PcOZ3dfiRWJss30rjk9+MBCI6zaUhCZhiNM9rFxnZ
JrohEa3iIyjZ2fRjkE38n65twDKRGfhNevty0qSp4FLHY+PeB1x5WpkQUb6qK7IZNOHrftxO5iI2
iqNGegkDjf/3x+HBEKIJVeSfBGcDSHlAaPTGeLf/npXam08W/rjrxRhsA6NB+ZsLSNZFCc2A1MHQ
btGxIUHby6RuMFPM6xfCtqbPiP+weL0BAqvNaJzxMLJ7C9qdQfgTAJBRKZwjb+dKnxkTC+IjH7+J
uex2N+SLB8fEWvJfwa5rs0jKIMf8R3qAskK7tRuAIKKKeMVA0B0CQ9KW/eXz3pyfAuHrfOv7URFb
pvdHzcs8n9/vytbPDzskgT5llYI0TJLfwnX5EIyM6M4pZIm57tPr/BtngYGQwkXt3KMjn3Ml7Alb
d55SCxSInRFRnJvVl4xDh1SNHGuRegsHGEDzd6wwOu0ppX8/XCJ3II+m9T53ZBtFVrZsdN6SyQQr
5pd0+1p0N113SRRqd33YnUzsQae6NHpZ+g9tRy1NRgVrZ6tsnkhxt+kkRKxyszamnaCVoYmRKmbl
UoIXRLFdf8L48OnOS0a51bplr7Fsd81SXbbyMyxe2IOOpDuynCgygdldqkLSlmE3Vlb7m1K3DU3J
5dmng6qTVLOAOM6DBdoHmfFL9rYQSD68KuXuQxMtVAnIlihExi1ca8awXyluP7iNb8J8MWiDuuTd
svWFHT8cFWIGdKGrg0HoEJ+0/4/EvHCK0slzSB+ja2HFJkf5FL+O+u3AchWuykMgphJbHBXM9+Yv
5lCQJsEo12kfNz1x+ut6E/5Py/ikF/FprZXQYz4iweHXKTmVrTCAVF8LR/0KEM6KJFS8cRjJLVS5
HIcD7YtbUQNyn4Wp6XmLFk5DRB/ctK+78lVSwIc22R02/Kn7bHA7Wg0zkOvZCbzyHreQp+o9O8Y4
3AtOtnS2/8c9NnVwaFDTkKlkDg2OdWWKetZvR43dQqW57kRVIRiA8AN9iTCvIkrnga7qDR6/UAQB
sG1QJ6rooLK4HJeClDJxI0pECKG1/SEcoCEbfEMkXT5hFzJYtOD1SKOY8fOVmHtopyPpl6rij7DE
i2Zk4V5Q4NojkvODGrN68y+P6ZuL7yOVoYJL/T7UojWXVWKFvShysYufQ3k6IuFIX3Fnxy5hX4+0
3EJ4bdtxOv97WUBmimreL+FM1WuVqz+0g0wQP4S9JhfdxX+PgiafYxyBXnAaehon5b0Q+DH9r7OQ
t/vbKohtVJ99SW2SGoUW/zGVaW8+rs0VDwoLHwQMOt4KPixSM0SvhEne5Deaaw+Ry4b1T5NbIzq8
6aaDanwmzwTPivED957KsqkgCTu6G4TWsDeG9V54/VZSCmfXSucWCEeT5nUHtEwWmMTo+TDUAUoI
Ghu0QfaNyj9Gias+7G/ofHMI4YuLRuFUuC5b9Xf58EDkgOTvp9mF8MkFgr0LEg8iAwNB3vHWhCib
5i1Om4MVS/ipAzjXf90//RvfcU+UOxAuRQ4uPM9k/IZ6y7AdTIRERcUKVqr9qYtj2AoXwQA4h95/
rnsu9Yxqr1joZ/eYQyKGoUcGGw9HSex5+Z2/tWb+r8DCmp53DlNNmEuaeKvFA8CqhlzBocpH1GT5
4rkyLaQe2SSFkbdBnoHJzKf/kVkjtbZBpyACyHM0DxVvaxd9OcWFhxP+dtXJZDaOTFkzrZNV3PFT
sAH+AylMkuAT+Mjs0L5b+jek8VbWduH85g+ZGVgVxp9q/2JhpM2t4EmMub+Y5nIq+xqZiglXYBJ/
6FCRE9zh4SWgVOSZC4vAiI8lnV56bNW9gpRUvfIWjpD/1xVvvHecTzr4kyc6poZRykaheWwUN7DO
drUKAF1v8Vt1xCSGff0Kx1r25wiqZlJSNCsG5DpaQRvLv9g21uvKCF3BpblTC26F5x+2A+8+szIg
Dyh5QEiQBNyZiA27/nUvF90dV86NuQ62OaoZloYrUVBDptSpCH/fTUpHoqH8h5UcR085ddGYQaG/
44Lz7adDv3m5lDmQwD6ffTgbCJTvsiEJESwxt4k1geo96QEqxkX2D8hJwJmuWRHfKxDVlGvBar0S
LU2VJ8omT6sJb7EA9SWeZ5I6O1dt9gRD4C2FW/lInw20eKxc2iaxXrLFn9hBVw01D09rw4ChUkCj
67ZAkEdDfyUnjMl1kEEMBaqf5cvj/0rdERMrNFhqwy2CjkePNyw3KtltGIJ1ht0cdRTSeIJpLA6+
M8ZYys3XjFtSsE/6p2SrRARCTF8tvKp1KpvEkK0rT1Tp3bzvFgjOD2OVdrWR0cIEkTEj6/POOcq4
OUMGH+fSJiCH6YKyH2rwwdi9mw3Xo0LldyTaWlmhFuNCjGDePqLKFYfXR3cb+6Pw+udLli6ztRnB
nrL0ZfE6m4rKMS1Vrtl9LppqYrSw1uztUBaQBXDt/5RL+DFEt/6n4LlJ12wh/X/ab9T4FrFNtj2Q
8lxTtBUIprewTrfn/YLoj7bghpGcDAZ0hZOWPACuGg9SgcgqFz7ZLBm2wCu6TGUwPF1Mkmizkke5
Yy2PFx5tf9+4crE2hKJ73Nwq4ZaFqxM1CwuBw5P3wUvBjoPiPvhc+WtN0qGLiepETtZRTGZa+T7N
Cl7hph/AZcg7RVCuMB+VBS0z2yvG+6tPvWIyPkjpH21+vTLvBbUebDEtQsbLz6MCH0YLxlhg9x3C
2rGg4W+mS9lLJUqLX0uvkrTwUEXaL1h06WzAZC5OGxyInV4SJkS1DbGL3NtIAdtqD6ANJ+xYNVCI
FDHw8loYIIkRy1yPIyKo7hbUsgBK57KsXU0dYN9Y+kU9HQ1K62v7iX+GrJ4x9Nk/FXbGuDr9Gf12
D8CoFu8KNOhLhwIf1IR8M6m2SYDv3hNAtlJ1qY49zcN5f7MNLvceHHbJcLOD1cfAtxkUW/JKY4BC
dYdk/ajnb6NKKaeCiqa7a+0ydlHmxSQEnYqgHoqR2KY8kHvLr1sKRWIHB1EqmPomK4IiA8obXDt5
/Ms2cePHinIDphyCFwUjcHps/fNAHjPa0b0iKOata0lrfB9k1BUa+uCQsIgQ9nPOfbdBPh+JahOy
6WZ31u5HPZcEqpFz+fw39nMziKhRsTFNS5VmwxOIde84lWN4OQSLHXYLfsdnYHFNfg4F5giK+xMB
32BdIKHA5Pd5a0s6IELXp3GrbB4auRUrm6xnVXV3wZ0+tfH5rBgCl8w9zTnJ+WJjQ2DTCzWmR1kq
VsjV/LZ/erSlJqcD7ufuF4lkCTFF+7EFi/WI6fr3Vk4g8+dM5AGptSomg4bJnjBVXqNDwraZ4jXD
X3p4CSsC5olGzYe/J3wWGlH4ssaVqBIobbuKTmpq+O6XY3G66rbGvy1qsJtaMzVuRD7V0Fu/wK8c
1iZNInVbSXI0m3qqrPB26DvVUy5xalOVYBdCB1O+caszriTXOC4d4YFyRFtO1JyWBy3CKHsR7OmA
ntoxQljoJQP0JK+aP6eJHjKeDLeQO0d5iFlozvvk2L0+kpIQN9oYwpnR1PnKlSHoL3OZXGFvvVhT
qh3JY/IPQxp9+vTy4ERGB3NDnt8aNwuARpfs6rSmAZeoXNIh5xN8MQZC3BPPnhofSMxxCECynmuM
iml95dUtwS17rHWyDttvBvX/yLMaKy7CgPKzCAqMsW5KrRNo5yf+xoZt8xwC9+mvcCLCFfJmvhRk
kJW9hndTx99PJ32NROH01UluBlKXsRZFSDtBOamC7UGMrab6jnETWLJ82stolIT2c/T/dYw9uLOJ
oXfKEi7wGZHZc9eWGM4FGiXvMesHuC18bq5jsX/f+AYLdwED7ywcsPFiXU0ROOlrrn6cM9aWdntG
AFqOUtSMTo4B26uf9J9LIjsf3sGcLMqhA5G4RrR35a3Fh1XR/plrmcPxC7Av9WCPN/PPbIvz9LZr
r4wI+43meJroRdhj1VMCv4YQzY2Hi+sddWBhfSM1AVLjeGnSxILGiVm1M17rOAJVBbPsJC0ETsFQ
t3KN550yOShNZ+6YrhIUqFaPctytbZhuzKWdJgfMl4T2uwaT7I0D6aXnlbPGfzrnMMv5Wsg5JHxi
IqlPX0aZ3cgI3j8P99QP/IJ4MCU71JV/yZm8dbKlrdVtasljJ1Y27ifLpum6LowfcUCmMdBoDMQC
duttadK7bZGQmI8/PnsItIfh+Ds2QKl1J5ww4tCKznJU3R56lFaH7CGZl3DK7DpiYC/QwhyuYu9F
3B8fWXsPySG2tHTDUw+bval+2sFMvWE+aQzqzFiJuNNfOozP83QZ8tzNRauLfUrnlBUDejRuXx+P
7ul3NdkBl1rEsIzJLPn3gK8mXSqUx14yd7e7RgzAKdcoXRhow+ngStB5jqYlod16GcDXHu5WUf9i
2CfkwUXurtMjmP5CC6jHnvzMYrBWrUx4ZBK344d4aKD9gSpTU1IMXJgsAnGgZpBeCi0hxk6k1vDu
BYlAhOMFL0E1anobwsWrJX6vbJZMNZqeEptoyiwXitSm7UP7gJTNbGxtaeS4QgkmVR2VyPIMKZWJ
nkOa3IsEwFrBG6+u06UPvYspS6DvIcbLHS0UcCaDTFgod3zUKswSDfQHEw/gsqdK0akzYLw7sXE6
VlXPwBDk/S640rqwFZxlHN9N/j4T1F3CvSFgkJM5Mldbplm2XRBr3CGnkqPPZuAixxKFoJu2ZbFI
mLhX93xv8IPsUsX5aP5ESYGl+hCVoFsEZeuOE9dJ9cI/J96MwojKgeMChSs2C8R5VcJMcX/acaoh
yMMI2aeB8Kx+gc356la64bzC9Bj1a/33YOdjAq7qXpgOzYgLDdpWLaw4oZ9BsAEyQ3DIA1xISrvq
YgeyQegvsun2k9cVJWJ4Qu6GwdlGZQ3JcZy0qXv8Kt44QKjiJ1vwEKRb047gFHhSDtoIlsf3KBuo
qsVqcEluVlNzeuhR6tGgHd9hF7PxhGsdGh2tptL4hn86seIm9BPD7QJUjYm3aPpRt2iJjUKLCQV5
nfUS85KpyCWrT5JTSXbT29610mXr06dmTV1gFPfelOR0pGzG9fIggm/LjmYp0EliNSL9JZJfdEDK
1e68z5Uv7xpwRCYzKQeAIHmhsp/nz1FvGMTg9TfUS8TUmr6V+odXjDnz0L4do8eylGw9bSJ67RJU
Op//PURho7Hyzydk6c+HZmgR+SXh/inOfzq4+GG/WYiASdkAM11wmAwfzHxUTqb4r35m+uKVCOkG
bLQxE7qimeTqaow4XUwcCoWXxuHapSeVQzG9aNHfrr+Qzb7VsyAmxKWsBhWx4r746uNZXUfmP+t1
bOIC9fl6SCFwDYRrCf83foRoRGxDwb2KIk/LbJgg1NPMGnGG40k5IgFKe5TdlMlujJ7oWoCgQtj4
mHAR1cNblEFemGzfXJrdEO+o9nYVf/bkW/lPJzJ3EuFStDvpsw3iIUfd/JK5ZlJefXVBg1vD8vFc
m4YR8IuwaAmbI8gVMPwe7wkECoHx+0X5cNoKZDKFrHr0RR6TvgZ21KPAJTjfH07OSIhyZjpPJp/d
uixa2Jy5HPzJ/l5JtQmWgUkU6EIskgqvJFBaTVBGfUNTEUax/w/BPH45BNvXzCP5ejH1/U3uoFAK
U+rCuM1MojRu9FZQrdzyJMdF7wF+3Mkku6qOKiemmrvJuPpvMatHqHtzuKUOjWE+dKM9OJJJ7RLh
SYMSSod2TlhnT8DtX0MIdjfVVKBGmnOLPjl6LF5wTV0bJm9az10Z8cUO+QlARrAvc6w15fUP0cNx
evz6l/Aa8pvYu1WsUH/g/VreoKKNwiFgTEWuGPPjSe5jsHmmTHRNGOIgL/SpSGAhIphjUttPpQx6
/zMdY9f4jVZ/WoVVNMeq4ppWtI6XUXyb1ktBcLaf2VdyCmfqgDUWIUcus8eKbnket2DvzgYHs8Ss
RQaa8CpdyZCdSyUDX1Jq2JZicbMEitZCGcX9O1/jEUurbuvTv2WU7x3eytl16HBzPyhOlSusx3X8
+CQmuaEXiAVb8wLvsWG4PrWWxvAx3FBMZkDeJNXgqUQh+x9YJxQ4Qt2JyFU+9Lj2riE4OJaShMbC
O5E44faRlrorV+HfQvrKq+7qP/ogMVK9utFjvvjJEyBwELdaCoclN2YsN+hS1bdgylcx7QRHn1aR
RWXAkxwETg00d1g4o8zlQP9Dbgu/R2GrHPmH0aQP2L5mRLkmwAH4/fLU3Rk+kEQe/hVKDuEd//Nb
wxeHun+Bf6M3x5wL0seNDP6uE7SyfQH/GpzuU07puoJvOjLmFoPrIBSUbNgXhAqxo0p077f78olv
uMfhGwqvQXBAIow10bi9EnQj8rFNBbun/0QNDFD0LeNPa3vZZ5ktuJHD7IcoV5X2UiKSC1sk9JQD
iCU/Bs08jAjmZmBRx1fKtcegR9Hp76j0Ut0t+P84Hc4YNXwitawJ8e7CVEGeoIazyQo++wrwpm3P
D6j/fGGpWYfnOy208uv6HrJy4GCHoKeDh+iSPYw09dPAL1IfbfCRbzGqvUVkXVcJRy+X7/pEEcjJ
1iwgi57hacoWIMrFmyoeeLH1FxpYo/x3xAg+A2LQn3Kif0SwWw2vjhWcL0dzEzhWVIq1g9vRa9R7
Ad3Zrt6XO/wgbt4lXzHmLXtp3SCQNf3pb1ov5f/II5V5Kzbr1KEbaj7J/xGEL3127YUZ6C8xBtI0
qm6yIayUEV+5kCARm2Ejj5ppFCwtd9sJFKTKyEGH/589ktnpIHT6F63zaBmHEb4MljQRzhpmzfbj
1inM0/ZSxDUjyMkw/RThQoBsfGJ2tqBtCSNnjwk3+v4Qv5/mps+ULRod75rAvpnwnAp/xTfZQcC4
s4Nu3edvjlyqmy30kEF3Dpz1VhE0zZCYpW+wEszEfEUMFr3JenNiHu0TpUlKrBNL2tenYOS5WckN
K9kixWbMO9vSbbtauSebIFHGPejjXJn6blln/3+5nXwyy/RNe3JlnTDBlZGme1aKR/Rrg0VNdbGJ
fkJO5+LinkvDjfbKnRwOebJQibslcUlBX3gL6HN1Ymuf+eVrF3NOmfIrTaug1Vo9XueNgTvEmtyF
nm1N+dAbq+oWpxJVUbasgaavAtf56wX7S8+ju+gVeVpzEONVJZW06WjtLHqGGZi+6k/Wn/Vq/fsV
IVraaAVp94QZqnISL06Hv+1dy5DzNNcCQ/ePTDTvjzabLDw1CO06R8uIib1P8HO6wudwpIuqd9K9
rbIs8sE9PLfE41v6/IBXUm4WQhh5zDiqQ3SMS9L2ZQqFAGDYU8q0oJqYIDh6zi1L0i9PvENXFZxz
sHSLcxgC1kx0WrEL8bGv519qXMFMRO6ukAaYfNFit/0W7PmQh78SKScz0cd5e4DMyvE47wwnLbrY
e7OAYDZ8tJLf9S3n0OWrFuwPM++7hz8xU24dTM7emz9AUVRutgUWraagd3anpPX5kPSinkS3nM/h
Mg8S2OJXGO09YYikOkwEKEIy60UWiEQ98DDeqgvOplnubXKpo/z0vvzEfQfoSrG8cn+iVuN8ERyB
w39RD0eamppyN0D8Y6kWzpNWAvjz1VEAmRt3XOxK46f+axcVydYeJEotTSwtXuFe4PV50nFhIDBU
jOJzoMmhGW1YYloyFlEwlnfxq0CyJ3zyu8WVNTjXVcN2RazzHoBjaZQ22Ld8RwVPf/V89pKkMsOv
dvoz4e8S3tWczU2LrumNYkKeEGcwkD1rQ5wIA3XUxayWvN6AOfp8awJuXYtpk4Vy2RxjEqF8wVvl
IK5DitT/OPbDHisK9kfZHp8cGGqTXJ/ayrwQMY9y7MM1HYqEE4ORyu+ZsMdd64zbCeJmEPghWmMa
kpeNMU0k80AiNuc9vaP2Fw69d/XKOHEThx00oKBHieqApKE5tpe9vXCWvFk4+pIXNSEr23Xl0jJH
IyAoEpmVPSa0QXq+UIq9tZVb/by3NpcA+LmhRy05AtxHkvRuReecppUPMZjn0gdQHg/O4TvlMmXc
cdcJABEmRMxJtFeUwADKxTuXIuo1xs2QhVdRxtOIaD1+iuEUqw/2NC7N+N98VjQfwHLsTvzDZL7L
jCeVS3upLGCxpQFtgvfe7qQJXIdTBFIkdfKgr0BVbVfiSFaQY/I7l2/IieRmSoBKyns0+S4Ng2Dn
sfbG1nqMxxJ3rI/TSXoOPe4H8Sa7yCVb+BJ2uIPwrIIPx2aKspBEdyy2au/XT2qu3rfanZgwiXYv
O24elVY/o/EG6YgiMtrEC/IB10A7nh/sTEO5qv72V73pHqp6ubtv6L9uumn4MQ7RJB1RTdA5Ha5I
9kuMD/+6pg1A6bsZpGQiwEjwImHSwlntrLj7O7X7o+9lzk3y4y1TbHxMYOCjP0pOq81pZwgVlK2N
xUc/0EGmyaetwTGcM/qUwmdpk+f1I+UKftEPitNkw9hYo7tAH1nTTltD0UMzYg8xEfiyc1CRex6p
GoUI9cfe+YH+Rd3dO2KN135DF9G4csRHvaI4zWyP8VznFp9eVNWxl2CA4bZkV15ksXBhpDbT4Gja
6q9L5P17yF2S3eqs8Aa11Qp1sRDaT5JX8fdcMI2prG1xbAXX549E2F9jTqeugW3E6qD40AOKKYhv
N8mRmkmdmpqHW2fZn9qx+M3JkNh9/GKCY546arlMd+mjS27ix2LrQf3b2Dt80Enrm0pxtUShTESo
c2C7keDStPEGPpLFXZuT1xTWJR6G10xy5nSvgEb+IDhpfk41ZWdjV3Z+/a2BFUjg6HLLPZdv5DWK
diaZmh2zywQY38i3zO24eRDI4boCBFu7b/kC3lJhmrsHfpgAB9Ix9Bry/R5QNu4nEPUwZCBZ2M5E
RBfRkVSkk8nLL1IQuB6xYuCo3TWcfiRh33ZIh9VE6RoBD+IK4vqQBn9kuA1mqNz6qfizKCtkeXv5
YwTpwnDOLBrCE7+bb/4QU1gSwVXPGZXqpEKdKV7DndhB0yLOrbHScY9z+RdbLUWDv6uB/+5BuKhO
23010eiYCXtaVmeep2xxCz3HqKwBnoHnYsueFVXYohiFTRET+qcruuxxzB5DtVlvgv2hPD5O7Yfs
5oOehgl+cODAuWoqAYK3w0b8OXyaH97N+UV1apFnTLaM2iqSW/4+j/CJc2Tlhhq8o0V1FHaa2Q9B
WphekBW7acZ0zvbfB1/0KQ7pacnRnr9FtTEwJx8LJm1/crXrGOT1ZExvhzgH7Yf9qq4hwPzbC5OE
J21HmlAYYZEAFKi+fU6tNOQAga4i02Tk9/elSt6U1u1g8p4aOpbfPxHamwNS3dsv7p0EYb4XSSo7
x4fLdmTtfxw9ckRPdJO4eHT5+ETxLHPkzCSvgjif01a/UsN79YNDcG6hwWKv5GFsFNfnA8y/lkob
/Nz0Sfzu7qyGBqGyn4C+ShcQwUDZYmsWsA/z3XmCA6wMwMHnM5USXa82LAWLSCHPjOBXFFXHDScU
5MDCXFfap0tK95bXUlC2608q2M44JAwjJjWTf5aX6Lb7lo/Ci08vpbEymcPELwSpcWQ/6TY6Hlvg
9VW/lDwsIObzW1dy8peLK45KXzWiv+B5AO0YfzLBswFLQrl0M54pFpwiEqqHp79HdRzuWn05XvvW
AZu5MUolRzZ7wGJOeNEvcI77EbyI++pS2/duUuP8fE0WrkY2tWUKm8MG7ExXzwIJohP+haw5Kf0d
Xyj1Pkm2R1HF/iTmLqenqa73xsZQ1lJjc2MKWwtJOzR82TPVFyXHnxN/yydi9+e2yW3iNjESjTef
pdEODVEBOWpIy8qcJXn74tG790PUT8ZwarjtkVW9Lk0e/7TJCRSFbY4t4o1xXwipzTmyy0COJoDU
0PWMdFTuOWKyCEe+HU7ZQvVukXUzencpLSdAuHvBd7jylp+/jY89GiRuBAcet9s5k09rCyUHL6YG
7zvDvm6mlpZ+Xckfm5F21d0jIh+wOTzzZc8dCMogxUGVR1clAAElshRas6N9R2OoM/LfM8cB6y3o
r4sKqBHFMkIrk6m1reVOSIxzGuo97vGq4rHeZjW51pf+3p6j6khBsCrmFY68JtUMEznVbaK4+h2m
4RwFFYg9Dw50i5Qt7eIr+BQUSIaAlGrtgYQk3S488RBb8G+qzrZo5RkX5JIJi2h0P3T7ReceQ7GU
EYdDaDu1OkZxbuyfV+2WT9AKB1zob4RR9s/tPdIqG72P5i71fkWQs6YFZRqs1KabXqvMMnSEN6nT
oGfi91bPg7npl83gL/h7eZ2JFbo99277OjcioQfP88tErzJBw30dcVV32+FSKQl1kdTnAflN0U6a
sgVRQ/M5PxHDa+ewk8GtBf28ILvoq1pP2rSkx4TRHG/DKjFrmUXwcWMmRVf4NZBn6TS7OomFuaC6
zsw8xvsjJcvd2FEdKtg26Kqa+U1hI77opLUCBRa1b0t6tM7D/lF/siMugthR4gmHlOIANijT7Eip
RYycAo0fOaUMvOLizgYfJ7ZgqzFVEOoe80TCaU6Y+eVSe1ZZN/mnB4HRq7Q7HmbR86YgRaY5nmLn
wksJZBEiPDUcNkQMRJVnCaHRDd43pqTODLZjruQTnTKSLmk/Kp7Tfbr9a0hRsqzs2Yb6fd4qobuc
lEv+RiDxeFu97eaKvMf5CA2Yg3HkmSlY1E9t4RE79xAuNZeUqEzTVbzDDcujX+g68qU9R2S9AdgL
bH91HYsZ+ygR7SUeMIJxY8jpxprpCA2zmK2d6lF8b+dtni95v/zyowdLopG7Qi1j/j3Nv1LgZEv3
+rMks+T9Wz8OI9K1iOKFrauHZ/KoLgCOmFnSIun9rI3WERSkX6rop+jg0WT9Aex7xy2dCcAol5zT
b30dfQMh0EnOGENEL3HE5e8qVbQk4SKYwjr9EO9ByJoGD2l/8WJVJ6Pk2evsSY6E3E9Ci/fAbmsL
6hRQUN5Xqh4Iil0bUoN/shqYu/IjIDtGVgeT4R8AdFxgWxVnOt4OCBCtOJfJ7Ycecj1M4yq8zK9Z
PAC2xJ3s/qJm8vBsP2tl8X4bgEf4ZzSjW3bv4no4kDEr48ruG6rOcun1+QX98PRGSUGkXi6wzGp2
kWxnoECqrW0dv7Ic8xOuvTIajcb9UcYTspoqk2j17s5RImnihJRv8YUovHPM5kj+XGuLu+J0wJ+p
0vImGpsdAv23n6OdxKbxHzOAcwzi4v7dCVrJpbH7Q3pNehed1tBej0t8WIWx8ZSZs52gjslLdM2t
+6ShTwNhUv7CypCanL9P+Lj8V9nezQCDdcdCWxp4QVkLTcuEE7DEGEYYofaMvjiwpUwpl8KjF7G4
Y727y6DcNXZSz72UOvy1fvCN1y9szNL73dVm3e9G0mKJVnNrF9ve+XawfF4OFR7HioJ1pxE1OSbJ
V3Ts4plW98YpT/TZHZyW9wz8664dP8uA06jl116vR3wco5dwbetFr91DHNXSUjeTGrz9AvqHawx/
24/aYCaDNBKxHU45sAY38FBWW3L4pXJ5bbbk+4qK+3cD7uC/QDjPGAdsaHDfvp2Ph6qPozWAcv+w
tdTONtHShNFuAUa8oBFmneReLBNmkyywOHPDdRQ8rj0dgApjV9kYjXpUVBVMS/BSyZU6gDMg0+7o
VN1AmsHkVVPXIuPydToznD8Kg9k39npeBkrKZ6lVBsJBHs1Fw5GsFj/Q7uPvz6zDQxthhTYHxed7
SEdcmJ+SNKQGvDH+jkxsF+UM4aLcpTzlaD1yKIdOdUTOs69Py+PqBUKYAy2/76gxwTq4bPIdNO0u
9TdWirjJC4jHJxSrQHx3lGlduAPVTXlHWYq+Ks5VOJDChKtb+kBws2ByeDhtDMuY7e3yoaebX78x
trYLlBiAWpsh70DzYW0bhuscsjN48Tp7LFesQBmFIpBu1eA0EyB4oqiFnvFOyd8PIUA/x3Kri1L/
VNP5UJuwvg/7MWxn7EI3npSlW+Vxdqf/IdL35ldoCoBMgLaZpxtyiCCmkPuxGGCMQyAzZ3cJww7W
T81zanDSh0kS0shWnVSuujq5Ui1E5STmkGMVU8FC7NVGtZYS7l1iMT93RREJutRFJEQiIvSmSTTD
5X/IAgM0Mmjnqq1MNvfPJ6cIPpymL/Ue0SoJUGp9sgDFDYr+NZGMQBYGqV7BCDdIZFIHtU/Zc0G5
xqG/Vd8QzanIw8qzDO8yu2euxANHBhYJ2Y/0wbflcC8OEl9asQxqr7zgDWvkusc3rsiTWhxuxq+O
V9NpYQVu0VQl53it9RvsbOx3jWREeLujICZIdwUQ6Ekhwu6ySQei81XA4fPckzLGrlnH2eHd3pP3
/IMxQDONGyqP1vt6jX4XzQnWDWnoNC0GuEy7ziHD5y3VPpNBYlgLsDZzB7fkpmnGYi49MdtlS/tW
o9YDR0Bs5dSS6Y0BLt0yxIEreaHPIQ6XPJ0pC5yM28gS/S2ritdAda+HRgfjuJRm49MFPXuISGP6
rVutV5W9aD543Yq6nGNNA9s6QaIWIcfQBpn3RgTjwltL7gaIBhEDwtRLxyf2YUvIdPlGD+aBeDa3
hgI7TD38r1o5v5mYCs6KbS7XW6s5VgdQ66hCXwsjbtG0vFVi8so9TnB8UO78XtZIRms9CT9nbH5y
nfRc9weiO1UiY7DXe6/+Aruaf3M7AtGHHg4VwoSp6lBOpV2tba8P/U0J80LSPxt/0Ycsa7B1H5kh
ULqXbdhRQB2Wg5ycTGoywGr4r87UBHQPN5w77vkXeIr8aIFRqs0/jvaJIqFHJdRMMvt7lHGYnR8P
z3137dRpglq7T2d1YDkELTPjtwVtcjADw+1cxD5RqvY4Dz9EFd4X6TNRlrvrRHkMz+w0zzq3DfEA
L+8YDvyedKldOSKpUzAiilhJcGeeJU3n8rzX11s6djxO4mh0D7frUeMm6RCAFoJjuPVvklSblerc
AFuuT5OTNs1h8Byrx7DI/y2LRzoOU+oCXVhUs4uBoNgHsX+ASNx8nDD2+J8UqkyTcMeu7m2HgbBr
P8JeufseJ99qtO1tzzRLSTLpoLe4dWhnNwG6J63KFIS/dAZpg0llOxZk+zy71qewHVm2CAOCBegu
o0r4XNw6e1t81gBCJFETVO8xZj7S3ZhWWdZIgVnawpcqJIZdgCqQTje7yuq8LgRsSDS2J4BX/1UK
j1KPi4+UhBsvstU3MA1+qnzvH1e2CNMMN966EUqfdWWZCD24JWunCw+sdjNmb52+8LvkYTilGWZS
v0hlAgcxg7MIDZuvbttjMYHM2uYDJLULg+YFmQsFQZvfR3DaYrczRVLHT8hd+Uf7MqrV9wnNDtcZ
1KgJJGyVEaj9LvpUUoQkxgH8hH+LGkmb2b0PwYICxy2Mat9f0DmA+QG9cnzgpRxJCKGjNc6p5WSr
mC5ZOBkX3WUrNwRO4mT6qOdT9br+cg9feNQLVwTJT89aeL6TuzeUUnK0HAXv0Qu5I7D8vmJN3sa4
LCiHXJLhP+iz6tgmO1lNC62xxiUGt46cjv/42PDV/GM/9MWUqIJJZY3mlV1gJAziXtx1cocngLbq
yN9nP1Tm5d1SfRkGDSfNOpehRdS1vD5NEKdd3Qz7vi6oYxVwrxx2L8RBZtY5AzGCEAns0IJpwShx
tS2l1OIl3KeQdvdNgmN5LnK3Zc5MiFIiH3L7c8EKzOCJuSlmziqwS01vH0x6tua8elrakPkTQZpS
tcgb8BPa5Pekq7qtLKV9FaAo+KLFp3dsH9ntCkREIEh8Sg3OXH6t4AVgi3fHZ3MY0IkJLFnlvzTB
MT7XEIPdabqh99ImZOQWSq82prNy6rA8OwMrttJjyMIuIog3Ragbr3ZWur+6O1HSJyGFjjy3e970
X6zP3UV6ZSKN9Uis1InCMS2woffOr+pMqjmYU5/qqeFnrXfzRfpuPi36JEM22v3h/QoOVsG0wYLc
QCe69xqksH7l06DDyHEFuI0uDYjraXBtxhfKRtM/wdssnb+2esg4GtziEixKOt1NURAdg/aLyoro
AT96KxSnNuZIwdFBAOfI+WzCRbhBj8OX+DOByv6F+D1Y/FRT99ZQ7ZuQMZbk8KBKVnsHrf9hD2fd
Jd/gDAjeSgciRQmzmst+tex3EwgnrlstORTAqEidHlACf8QYrnZ2EnrSyo5YlKIgiosUuzuEl/Ue
DQnqKa7eJ6Y/3AZtHqmTwhcqNcpFG9wEuXM+oL1gtRRBAIe8nw8UbI/u/EEC8jBEPBfKapMByb4j
Jd7HnbSW3ziDoAeidM8Yl5OZaMqOehjQunlSw7aEoI9N7a/WDd/N4KeJjdMOuYQjV3ZkAM9zUKRG
88fD6Xp0IKzW5q8eQeQRVnKy/qpn1beJFohZaKCLCAvc3Z3GtgTt3V6DButtWhTiaIGPoliuEvYZ
zgODLKms1iVN6axlbn46tuzGc9nUciXjLvUAPnGV+ZMzJE5proVV+uBUD7wm2fn1DND3RkEw5v71
SUpQ9KUxUelNvZ3/FegC9bLZp2WvkNP2gHHBwE5Qki5OpDZ77vHRFo741FF7vZMdvCsQzDUCKYbZ
I1/668+zM2VbOmLpE2Pp64nwTbqnXQqWplwb7bHtXgSoWfPD2zZAewWEOvT9vI0Xic0uw2zd/ZxV
DNlxgb3daNJiSETqtvYrXKVFukwwxHlfHZrpjUwrZ7uajrivss3aDVF89o52TiG2yNAx8d2yJODw
Nus77IKuErLv36Pw0im08bJXxR0oQDGd+SpFHAVMNVBr7P9hqK+XB5Fj1t1iW2FXvEnRUTMY1qoz
MATcgHHvQqVpZ3EgR1Gjgslw8Ma6oiuFIECa0ckyFvd/gojyrQtaIYtT0JpuK/eavav38FKVSDGD
PlUPeC+463l/og5Kouh67YrEVApmqIV5tt1k0wDBWQ2RUmxr7OSLb7amD2ct8nfgDs1N+IGH8sOU
6J8jjRMZOdqf0gDPuvHS9uurp7SXrtro/OILICQr2nmsG+GVdyqmATdsb+w2N0v7/gCZtxnRJtNm
BfULZsyfXI9u+JmMwMhOkXxMa1ABx7Bg4hf86fX6fjogSxAnqz8ZAL+EkRbKtaTx05RyZX5FuQV2
wkZUfsPSmDO/jGn4L7S8b70oR1UeaoQWctqviVu2RHoAF/gr7R6RTsL0WTu73d/M+oALdOeKRa1Q
kQ1hgM7sOc1RNjA/SQ3rnXfUqDJiFhUg26mkAIDMVECbz5bis/OzpAVaifHlMBc1GfpxpdAnOt7F
egui65K7Y4CPNUroJtG5VtvCn0x8TsVx0FMi81xt0cj9cH961WY9Hyc1f6cuTO++PM93LvXb4XN4
xjTOVTDXhA5huNdjd9iSCRBQ/fScJpJe1n0lFWtr/EAFTOYlKAKeWffUH16eZqPBYD9pyUOV4esN
krWqEarPaSdFGkPk4aGe67SYhRYi2/y0TBT40NFdZcPlFjLiesTiwd4npy8OYyjfKnKfG36rWYC/
WEJpUr1FCj0PTcVEFCA+jwEnUjYaT19wjNfEO7pbX4ytCsoL9kKEvIyvSzOQmB5FgVGjb0o37mgU
HkBgekw/H1YeaMQ+Tvc7PPF9XassfDIx+qiYZd73bckoKW+LS9pnkerP6R6Vp98eONvd5ZGRiZW8
KD0Z0WRwwq3cC+kQ8GRKxZTd0NHKneQmDDzaiDSd5qJoxpFZfSpLn20JicrnZ/J1X6x9yHF627zz
hxsMsN1Yh2KhS11EgGz/9qp5L4Q++aOUOF3ho426SR4Tb4EXRldaTFLHdI6jszI+s61RL/2ZGpSF
xgQxJ5kWB+gNS9yinWARr76+nVATEweIx9ZrgDiZArep1MWQ/McF447AyZCqmq6e+8EH8N2rEDrh
BDzElcvI4X2yVDrKWynidnksk2L0dcADQTdmzc03NUA1ZWoFkI1JUmFtTd53Tj7Z95LOb5hYZ4I4
uq1bWdCEHa3mhQfAsr6CFBb/pLw/iSxlRhCjLm8udaFeWjapwuggTUgs49w2BO3X1mtiqThW4gcw
kdXeugXbhOUvFtozOpQtfUAw5Iex8Ev6+IF+Kj044/L5G1X5NiuV+m3Xt25YxR9tsmUEx0k8z3dW
wGstKMMZ71j85+1tmesUb7I60r9zVxWPK3HtvOqvsg9I0jQTiPm/KBddCgF3ptWbBhzCjxt5TYTJ
QazQNUyNFZzu3B310qPxOyVwoFY5fNwL6fyLt0y9KKvqxSaUJa+xhQThJDUOaFa+HaDg9KXPRqZV
LyekL48xjPSySy+OAM6AM3eikcfB1R5iKDl6pfsPnxuR3fSIpnvcEVoZmiIvcprqqvXDoZMTkrdr
KRnMr2WuPxfnXueqRM9U4YYWoZoYGWVVoMaUx2nMqDLorG5NDQxUgvXvU0vnIrDU54hO/mTP3n/s
88BIJjY+pE5DUW3j1F1w5cNvh6dg0v5QJthKRiM0Ei3kiKjt27jsoMcmlBu5s5OOHwpLbaOAXFiL
TmQeqxu7JYcra4wm58POjkR6nfvMwgw3KDubRjE+T0iL6qiS8eUEbLv+7oUGJ7SnL24Xgmq4hNEn
m9+Ox3pTOAhthw7blGBjDLkEwh2W/NfFSzHcLjKQ8JT3aCdKioJZ0htlymkPOQyiffgGgZX/NcNK
Ul+p/uWW6qbmZNCYeb+YSNYvlymT8FNqjxqb/2WUM4F7fD2tH4uONtSnDVdP/ZOAJZ6S1piqNu8y
ysDfHVjmvzhTK2zxLQdZ+Ru1kYChoSxEXLocsbRna62K32iPfRhF/Seg0GwQ8Dyj7sBftxv6l64v
tdg1mCXx1CLgvhMqgD60c0nZa3LKNcDr9RhttsZvdgJJaOCc4AOHWmqSDWUc8C+mmEhHfAvvLAVE
gKf/jzssIkWaqBmzAEZMAqF8hx5UNKEOAp3pK3w6KET/PcFqdwxL8TFB7B4NMpVrrhLI6qkhUpqW
eWvT9CItR/eR+2izb167Y6eYcSolsnBO/J2bzHTTsBasCyP7PhtUGwUQoXt8E0Y/BqSMxxnaJIJu
bQ3xIzbyBnjZUJ25MvIbik/v0aSQqVQGJGynpV8OSl8YaXOYlhkoJ858946QTrgKgofDBQ+SZfxq
dGqj38qtLSXdyfuhC/E8Sqa6P1f7IX2k/HcKKiProo9tgPMapLrF7DI3f4a+SRuT3+mIxULAFWjT
51w5nfY0+q7IVkhG8VbB9j6KDFIshF8x8G9QOSCXbSM0sCD9o3vPm0J6a+X/Jgff/uNsgDqIOiPr
hXq66IIQIHbGP4KqW4R4RpfG3hZ/yGEkQX3HsJC4DXkVibnTgK/u3QCXzmobWGBmbW/spri1Gdyh
dbhr/5OPYUVdhDvSVWeqIfrfOK94ubsH5jZbvyCWKnD1XTv3tHso0vU7eb/b+R+0PLQG9SLhWTHE
vcCkcK4GyWM9pf2K0Oxzy4Lvm2SoMf0EClT0TGSMO4Zc/1XvUGLIcUCLQE0I1PucpO2+7bBbmdH+
TM6n1EJg7MWWkbathqlnzSZ87cZuHI4CEXsPKN4tMyhz1jUfNfb2kgoqpDBEm4OvCHLof65dBMt4
kztlMv/XlwObdW5ruwLfg7FpcQwe7RUmxPov06y0qEb+ajvJpaXpczzeqi5r4Yb/W3g/dxsLbiRq
O2TVK4OZjmwdCls8lC/nULopLlkg/s5zhoDIh5YJSBxm0aCNwWUgUP9xR+d/yKgMt/xyoiQEQ4LR
AdAaszYx4ec35nEieEW7SRVpdx/0eAs0AM+HPPw+xOspyd8ncDSSEBRyFsD2KkJSUDQGzIOa2Ywd
q+5OHU0iy41balMMdKn2jYZpr4xno/jhSBJDtrW+kAmoSmQ/oRcPV9ZuqZlYcAH6T+rRBn2Cf4pm
/ULrn72JwvYwPi1mvnUNxM5vLlt7AosLqpph/LgYo8RMbgfv7g71jFqLPkaIKC7OXilZq4aDAqXY
ms/oPwikWCb1WQh0QFHgeqFa76kBu0CxSWPDpvZ17aN94XUWKFipZg57DRKlhu3U2Mce92tdaHj9
06Ypv0dtUqiMJJhFgjEgCPVUXp/OiLI3v7PUZexA5sXTcnKjzfpVMtUfDvLS+3HKBy2uWjcADbSM
8wDt5Sv/4/hT5Vi5uM6tuOGUcrpwpTsOdB7LeEz5HT3SApwpVqvNPTd4zY1DnnE0Vwo4LywlKE3d
AVKkL7YRRxfmFbKEGoTOdgzyKkzP8iOU44TZR6Okn/4+qzeArQdGreSJngJ4IbmpuEWTxRMXnPwV
ttnV62bwicJe5iUuAHB1wXtC8HRZJ04/Ulu6OGQUfxjc2Sjel2jkYXI+m86DjCQ9VZ7KU1SmY/W0
uioWI0//ZSoeg+YBvfo8f7UUboErFRohEpPw7b6Jd0Kfnle4ANKKr+K/j0J8ZduEyuekKfiYoX5n
+jgM8IvMGWxXwZVyTPgAXKTxa0nqwJGtz5qHcjj3hDeyw5TZg9hKPLiTl4/jHxw0vOrzbix02VmD
Lu9gzzEkHsV3GgbFiswRmCvtp8V34482j1nbEGl/pTyY9SRtjVWCqMnsNuccDCgPxxc31ZW66h+K
rn02BYquVVMWcveFrcjdNrp6E474Il9R+WP6xcXwrbTKAz3eTO5/mSIXPGE9vi8mPRNuAFsHFNQ2
UD9zm3vSsdg3E7M5le5B26Qn424LZKADaptvToOvIvUYD2H7cGqABWwXO8i2Tfo91OPYDO/awGsY
K+sWp/HprEEK1YdxHVoLafikUfqsk8ZAqFpa99tg/i1uFhWZsx9qiqsQBMn6zmprDShdRE3Q46Ta
8chIf64lysxzyyuTV2TT2VQ+Pp004Sw0bO3jetUi/fxn7o3NYTjIOIby2qzd3mLyJFifbd8j9N8P
8lvYUGofAQswNIo1pjXf1HfhqHNTjsEqherDDVlyVa4iuH88WHi9Lk+f2i7I9g8ia6c+YgmnEgxJ
Uh8N2Uyha8jrSoSnUNafEPfRoTCV70irL1NkX5MhU0Kz2gLFXy3WMiZXHr8PL6DPL9V0KPXEwXL5
WE+qSXSmFokjXJUYo6tqmnktorpWZF8gc89u5f6CesunjgOPQrLtRAhfM8WWcbHvd2aV/WQsmoDs
HTDWVqc42tSq0RFJTVy123SxNBOgbO5ENlkdVr/ubAXgqyeK7TcYF3UN9X9ZNNS17Ls87zCc/+rw
URGQa9Eto0g65zhA0CGS4M+ISJw67OUr2wckZlKkM+krb8ilG4nKptLJma0mb+MdLFYn70vS+ckz
jf/T1Y8LNwCekcNCwV7JYJhEf16Lv+CRtLCUbyORj2ySjmUae4PHX0J0naa5W8pdbCf/mUulQx9N
WCAYEJUgvwlbffBgLlyRlFhk5nQeW++Mm6p0o6XQlSMoIHP2ZCYazDss7pI5b5ws3GB3Uih7FWwO
FzvIKay8iECrfDMAwDDCr6JB+NMas940rbQ8rs9zPPpzWDd8SqqnX1OTkZYyl9F1NdPQFDc1y/1E
fg3iQ8RUegVPY3U0Z4wrGE3FdK2e3Q/jCP7MGjZTWXV80kfpHq1BHH15a7Yz6MqBiRsT6lcIdBXt
dO9MSLBw+vi+KLRqdijNEYADNcrX3lcU1JraDPZX9MdsXo1R6z3q8pvnOI3vWCfUCb9U5GpJkbM5
WaNCak7IUfeRUEvxQrmRlgGAdQzY/qTovt5k0AQ0iMppJTDA1JSd0YmpSsahqxxLCgFJMYzYPx+h
MCp6RsM7dr7JgAN0po9Wr4f1GahsNfQbk9H8fmJvwF6GbwdK/qCmfSl1wEJgtw3KPDuz3OyKv9UK
qCOBRt6uBA0M0LD/6GqE684yHmp4SvoY6G3+FIooIMn5e9M4jNhCUm4wivba+NuTRD+OOhiGYreA
HVsQ77Bp3cROfx/F15JQnWMwIbv4MqnODjN5gUtUPLo4ODqccTl5+rJ0hTS/JHTZp1S0qqPE1QfW
0daaPzUCZJIvf91hkRllwji1LTdWXuZYd2O6x+edT4INJC9qkWNxPg93XRJA5VYk4/BRbscW/9hp
zYuGe01EeHvCV+/Vp/sq52T+b04tPepxJMQNvoF4y6yJKZaiLJl+VEPnSOEjRC0tJ2khLrfUVSWw
H+qMYzJsC7A810Is+h4J6mEItAaFfmIOt7w4HnLtgLQV5GYPX1pkveXDeJ290BGOzaoQ6wagEMre
EbZWJ1l8j5JmETfvlM04faNuYc3JipgSAY37KDbSArAfAVYccowszHw15pwU602rBtlbGrzU7g7o
r37m+MH/hzC3CqtFQnj1rtrfTd5oLri/SC24hqtFUmSfUNWi5IsPO+/ijiulla8RWHFsW6FqxZ5i
2x3YUYeZTXP3jAgmvn6NUuGUdktZIRFyz05D5HzOLCDpU4FSiV9u9kPKqgYJ25PZWKwzHDp8iIxS
quDoyUQ0TSuAcVLZp/SqrPyUZl12JGjW8pR8BEHYex9uC7IQe5qr7DJIRso/Qk+WfuIfa0E28P5R
tQdwqoi0UJlGhCoK8ec5NhsqvPaefgziPRL2U+hfxPT/XIO9gIOiPMeok/LJWw8g0ZrpGDKrvntr
/B0OywktfE4eJitDpnJ4L+CrAzUNgI50ZfuLaK0PZYcr8OniARC9IPHnvBeDo5/C1opygVf8Rzuk
bd1HEshXjoHdM2k11ZgHAF6zSl3VjT34/S3+tRyF62U81ygZ3qYi2/6av1+CHBOYPXN0xU4l6b4e
XtYT9IBErTRFFxOUQ+DTRZFw98WsxX9QmLzktW+umJwJmvvBqkBRrubzeFIkXRw27x5SDmd6mL7S
YnaNz9Zk3fMsXGvpozg1nNoOrgkwfsFMdPkXJ5JCXl+5Mak5FHglX54L/YNS6YJuCUZBJUONwpwT
wu5W8IjkCqk7Na2j6i93vd5NCLgzvwiK2tm3Cl99SFcRWiNIQmwwUVeOMWVyjWCf9IpM7l8LMckR
RUVVZKxn3KXA+HP3/HV6V6N49zOeA/mXmwun85ftRusCA0dDIUzn7R7/HknP1MjXUJhHX5ViDHD3
tJ2df2VADV6THAagdmqC5Y+6m7lIeSgwh9Nh86KifyrLj2BUsONHcrYqXpiL78PQWN+XKU3/1HuC
6GMCOqBvANDzH3My4s+naweVFVk1JxXjtsYqc7mbTi+XU1FEMYlX7OMgdkFk/V/sRjb1iijzJZes
3hmY4sEHAwwu0iJZrORFpuJJbrDB1vqjinCq6Q5bvBHRLJl+lbRyp8Gz1+YF/MRpi6RQ4K17+/GU
EqbyWgq8qQA1p7JKjkdxd5E9edQO9sFiPmWUGFur9saSWXtAiCaQE16comya6CkZAufy+BzMzZrX
hmjLnMGosoz9qCfuEnjm2blN2P0q1/sqnPP9xz93nrAxHwm4e/SNwcOWQy0XPV1X/UaM4ZtJ/16Z
HK9ka/Fx3SGtXDGswdlQSGoYVBQyPm1prf/FSe+Ajwc4hwCyJL0FVe9OcP5v407UJJrIIKvjjcMK
sSCCApSz9IvFOJhn6FEox6DkMe01DBbqVFe/4ieoWsbLOQGgx7DRQ49UjulSwWmAoXRlSr3pwbAN
ILaGTiNwpXeJj0hadbej6YUPwUi/JlgGoKlzwLyvkELtZHtS0wKSYKxwMtTcRxbC2PgYmnj6j8l2
iDnSFWTkjBh7YLYMvbzXoR/9GMhnFBNFEy6xYvCZsUg43C+8H/Sxe2BTcqfsclN1JCaWRgVfSVUx
mWzjpLBnW9kSzvP8Z03xUDRcbEuJ+qRUU8yCpk/2Hc0FDn403YNCSIvVN6f4rcgXwbWsdqUqB7o8
e0Mz4EV9O6T5hgPNe2L4sL2gPrICBsMYYqLBn8Oh/jkPoF7jrTlJhXTnoisE23obsEAZk4xUQh7z
JxMvodXHBjizMLLxed+oDV7BUsFKAgZXJQe10fo5ODIBePOKMhhM6JQME/wVpM2YYrG0N5BRUm9a
iuxSWf5SqjEBcKCVaFDNoZZrJrUBjfh18wlcQN/QXoKZKwKpgvqBMaAw0q8LDetAcZUuC69dUoTK
kwCVO+zTx7HWgqrn6j099aL5OvN5e3GNVwmNJ2FgnpXNNYvBWjISq35tEkFlZVOWc4lNnHuhXHOD
zcRQjzQeQ2nIdlxfYMXSZHcyvEfxt8/UW+RH4I91Pqvdg4I9lOi58S0Fu6kwpBe0voXTWZuSqDJU
gQO6RwA1jRKWoHZkf9RVKgujgPAZhHb1xKDc/BDUYFVIbWWxxHqySyeNWjx+hvoE7GIvRlmpyWz4
Qm3A+wPVPOYN7ZB0C28GthCfgiXI4y51lNOLIoXHwJLhC6H8BDOIcEoEW/aMu15l0dxVAvSperFx
0c/HX/oDLKdwhJOwOO5SEy0NRDnA44d+yFXUpX64cPChX5L0adGlBl3Kpu9/glxV0S+wZ8xCRqpP
yw2YueeYh7jG6Z9kNdVHa9ebT9doxsTUPdEq9C25K2fNsMX5PkztmGuOoBiJ93j6cVgLyyJ7Mzdk
2oYXNpilUN6kJhk918HNot2c7BzDHE7/V2DGfxA5J4ZYNudIoW7WBZODsMKvyOvpO+NM18D9NssS
xFnIKH3/8ba1i/VowuWQ788wfvCW72MZL7Lu8bu3YUXRoeuHPtx0wwBvZoq+zIwTUII56wnb1WGx
SxFW2RFNxgJYKC9c64NJ7mEcWeBUtpBIKQXJigGXbP+2796gFGM5pHt/DxDNtPDIFsc3S0YTPxB4
rz9egk+trCO89aFPUW7e8TREMVEAMbxp7uwkNGLKg5nu1QZMXqbwNLsm7qO+o1dtfGCGardc0nW/
KNBJ6VXj84CkfUfM6k30zFBGE5/Uz+69TnSPla8E1jKLx1GyAOu7Xw3y+w3r8NkXWxiSA0r0oUgm
n4IFiPSEC1XUef5PurReDjF2gKZZV1uoQY7i6oSR54RiZQhYrAqtc2cX/VaQ9l5OO0qHOLWibPIU
SH8AAn+JNfu09wN4bgwkb7TtqSyy8e2iRdXlISeWoWMM2A0HpE93hFOFl6QB1uBfsR7P6VtDfioF
w/03igNK0X2POE/M80TXNpUjuO+GSxC1cNS3GQSB5jbSJVts3KRk9xyeRQu7PHva5ovk5sGgSq4C
QnLSNvcv4TJm00oPfRe8aF1a6wr+WCmTRpLzi+b9VF9v56L+hytFKkXxPqSqbKC4Gwyus/LX29p1
XtyD7/C9vANqr8u0VyuBfr8foNjfrY6jY++JRmlYbqVw7nTNNlGjdWPSf41jkzgCtNZgS8nzlJmJ
PvSB6GXDzx6NcOEu9paY+r2h3EuBbR3WjEGNT2WQvSgKj23UlcD500DBXTFq5jv8lksvG4LHiPNu
Hjyok3Pt6DKiz3K1okscjBPnS9wCo1bvZ1gTY+3d+WvQ1LKrTouqARlcfeXU8Q6jPHH8cUMTlTGN
6zy4stdAaf4k80t23Dvs86xrb+xAzgcR4SEfRLpFVGlSbopZHK0YHjTDlsk/4N3KP2x9imGjF4iL
h/hRVb8QQg+HcdsqVJ63yeXXCY5gzSYMWaLPDL+6B5FIsV7OHkjKubiN4MwrKrSTGvfSGa8SaERo
yCP3jBHaNFel1vTRGGVDUOwHYI/DWERlXR7BdbAIv4LFXRcgv+KAQ9v0ja/yuMKkNY+MI5H1OwFB
YizNOelq2tm7j+3Ln2fSjSapLp16iQHYgdTqPOOTlcn8UaBQIaHv58dgbbQdGHB6rC/YPQKT8vo1
a8+Dcq3HdRFhD8/wcBDd4TeswmUZE9md9geb+DEeR05N++ADcrr35uRpn6XtrhWHBY7Nc7tCezu6
/ZZ6LqYnFSY/LjmcxjoijAP1fve5G6rYjdCK8CVEoJmQI1YCwSndI08e1FIZ3eRs/RXSLJVXd47q
84U6HwH6ilj7uPETDHQuTmEsJtw6c7oMKPzCYwRsjOnDOUSmpJr4eJVP94BPIPkcQNCF0p0XHZH4
XDME5urIOTmG0tlXA+on7nUmNyD2MlXeBZ3nu9naIKniHAJXe6S2BU92uWz7FlKcILNskHwl8ylH
BacvYpzAocLNuVGKaqJkaHYdUCXiczQ93bpn6nPENNlBB5ExboRsipkw+REtrGO1l0j96JHPqJJH
47T3t+FrBx1Ag3rVPb+Aqg/2MnCtdpMg0MAJQChZQsBU0dIkVdbuQIbmVSxHBfg6Y9QfIbQhTEyR
DeDmsm7FlMsKZfzJO46Rp2qhMTU8o1OwXea0dfO8wmu0d1VPaSJkbricVjSb7KuLG7xU94UmsVSD
lhUdGMfHNd80gYT7Ut4A9NMG5Q4D9mrDjAOe+LBW7pBmr7FzikXm+bhpVHFfuDHALSfaGEmFq2vJ
xZcIQn1LB9RnchaPbdfnZA+dwS0QN/skaU9xxRFbA2JIeDIGHL15FYS8Jz4CsKPAERb+6QVUmPMa
kTXT8dZPv8nYEAJ5ArWjR83bhTQkrA4oZRa4uhI/kdeONbgAPEvm1Aj8yf2w+ag3kOzbfUG4u/JD
SiVpiWbhC8378YE36cqa0Ox0nO0GsvLhdMheOMbt4WiNLauMJD3sJ2D7oIpdtAwxPbutp17I0KvM
8D6CRunxFM33hGxtvJpqZoUZcMH6DhWZsYP8UqcqZWopT0cd1Ws/Ggwl5LGF+aT267EVQc7CNk/Z
oI92UigofE09Oha7bxyZB2loFb66E/N2RGVmtZJ2TpoC3rXww3U7eOwNlj4Ut3SzpJYUet7PWMtC
mARro9qBiIiP7CadGvuBFyIogcS8yJHwMbfZRLCCvqDWWHmHXDm7Jb+FxCGgN0Yf+sEyK1JU4fsZ
nITCk9C/D91A2QRibQiNva6NJELU/MvfgS7uj59OPKk6Xq/nMTMF0JrHJvB1lpQKYrkeAyiQFtBm
3buK9rZSYmpQ9QwQI6J0kdcaJpzYxYb004LxwbhfhLpbU+hcTuscgZ+yhUOFAlVv8sAFgToEnSDW
OOmN3Ydt4fI70+HDi+uratJnj7+2SishfdfwljVUQz+I2CJ1RN5RjaWJkN2MsajCA/tatBVLm+Mi
cozx6i/XmVdl2XunvxVtCDYXUTeCal18cCVWVGehIv+39DHNGA1C9wol0mOMPpR8UKs2mmlfpePY
Tu/x+ElpEBsbunnNpID+krVtk28igW3Kc/rLmZZCKWJfILiUMHwXYgcKWCN+7YwwFLA1UjVaw9CK
4+PxAcKYS/3ZpOaP02lvMiKr2gNqh5opIDnV+o4wI+QE5a+t5LueG/maJmPRieMa
`protect end_protected
