-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ybptm3BcuFwRZai7Sqlx2TfDEIx6de71qflZ0H+djktcdXAtzMVXxmAz+J70vLTDRE7wcDmetDcN
n8/JxBfLspjyAouyjjEhZ3BQoKfBWTMWrz2Q7eL4WhwLyJwgw2uVX3v4W0Yu6rDOjuRAOCVwPAhV
vh4vIMzMI1juAsSHiKKfHs3kBKx7UJbO5bUafzGkd60TINu5BoW1fJUuNrSCAhff1pmYnOsOHCSo
tanfOoSpNycffDstO/1eh5SxA5L9QGFuBMNaK138C0jmZGCL4nlp9Dlt5gBxSDlrq2k1q1Bm0CCm
lo/Y7XRUOoJro+hQU8kIhdMQ/FZb35fEOK2TXA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24768)
`protect data_block
4YnkVpoaYXalSKwzUVvkgwNClYwbjubnTSbgjlX2QqwBvHfERzOtGMVaMdbDxZXH1/2OmApHYvs0
dngJcgjYsshbKy/HUE24+ZOCufv7cua6KG1lei3t176InhwFXUNEAW28+2tMrKN73aP2DUA4kOud
5IIeG+15k8rsuc9Xq+xl7Bwlo7JB3YfxkZt9tIHbJA/qgfib0nU5vzVlEv87LmM5rn079OiXXXKp
NOca/Iba8tvrn1BDwQ+Xm3eJV7i1/1GnTEldCr4DGMx6THSQ2Uvq09F1214+BTHtZWDa+bJFRvWI
KEUXgGJmashlbHwm/GezRCF5LOyLUawBJkZL3LLRNWsuham5zqMU59plR7M2LunrlLcMMM5CnrhG
mvQ0EhiiNb+QnsFTuFgH/qPBgHRvDD3onmsWh9ADpjKZ+x6w6kSDv2FBUk55/nnMEqAKzPtrFAyH
//0IJ/MLm5h3VsqjXOQrROQxrmb3/GBztGwgcZFuif+s6YUfs02too8LVyVMa7DLyH7n3ouNDIRO
Dsli337i3HVs7Py62ryo6L2Kh/Y+IZafRlBSZ/AjtSJRBp6Xhs/dkTAyqNWxxF4HvIqyM3MJe8dD
ey6iouJFb4O9u9u9XtOXbVlpWSTJX42el05pDHdaib2Jb385EljUABGxLgohsXU1JUtHu/8juIrn
6m+1bhb+IJgBI5AJxs7tOJGv4qe0HAC5mAkUbPtnmkzq7FESkVFrjPvYcZiUxubfinKXS2T72dfp
hWPkhJk7xW+YLLEZ50oCcP8IInlcy9zSJMfQ1u42a4reKiUyFbuDEU1x713C16CtTb86F5qje1mR
Yz9ird+Hf+m0JkDnoGU/XL+jpWxtkOlX/ah8Q3d8P/kocpd/YZjOCgxo+skL47sPhpYOexpj7K0q
80gjWRho7oRA/sYpCClxLDqwHgSvsOUjF+UNwUzlr33Q6OE2nzEDWbSN9k0XaFs3CKP9OQggsUre
yLA0f5TGLWSkGjybLDJCAyOwZUrlCzNizD09B1xxIcQVs0mgNx9qma3t4WXfCg1FvjL+ztijkhfM
tuW/95+ssGsvDIbYsuWXy+FCIkBqzY2tATsLK+f72xuaGIDyRLwDjwv3J2S3csC7wy6GvAhIu1WH
bwYeblluiNMTPVROl7lMQjXXLkgOwEBXyQFLBw+a+tV0Bmjmx4A9czfJPe1K75M+vMFSuGuLEGNA
/ZSGCgtX9rpECC2BSrPiGhu6PST0MydE0McSYAuTwg6q0DcgBXg/wr68fjOCa8hl571WLA6563xT
hgdQ5tPbkk5/VerQB6pTciadkL9MNgFYViqbcdTadccW3rALkryrMay3VEXIDlwYO5qNasGol8Kz
/+omvYfFAFKlNW7jazFbSau+6VKVxa9OpW6t1CmOGRsfYabDb45x80BEaVR9XDd2EYaBjA0VH78F
pLPGa4IEFn8FMcnzxvswU59oNEpf5UmLN1cm+gSM4EwiwRjPWet+iCcB4WXFzRWNb/VzO/CSyplk
b6uZlb2nNvZsD7HZtfdMqP1kxn4Kd1yTS4xfv2jGKEyCnJA9fEvRY00FTC2in5DngB73baLqq+kB
a6UMKk9LH5U4wmIQDi4HPx+TRFAXSJqGElsc/wWp0wCUp5L/EmnEPsYAtw+nVmDKrXF8SHoNa5+o
Wv0OasBP46yP3dqVAjyw/M28WzEoaeJAp4WfyMUZvbNCv7VMUrMpDYb1QgPQPNeWQxq99F8xaXPd
X/umXpmIElzxi//eQYHFwanA8J6bS/rUltmyNKibuj0UfQ5S7yJvAyZvNXhpxTUxb2BvvIj1rgrJ
opRf2ia8CKgfKWrrT0oQ/lMLHsUj68Ug6HU20DZfUxCmUKryCasGAidsPHTyAaSPLYZNSOInljG/
lrdq4YTZKoX/9B/fDjc1eElF0CKmnoDFZlSOKpUsq0OlNXnWa/tyXh9lNI4U9nhkcCgoT15Mvtt6
SO/7YQV3HEQ6sFsVTl4hJ5fwxVoaWNiWysi/lkRm2LlNgP2/9Jnx7dbq/++LHZGEikuyTtRGsmzI
cZI+yEXqOSL7L/LxVxg035xJ/TQEzJBj+JVs+S6VsfrvqJ6hU6QzTZCpiStdTF/GBc2Zg7Wcq8hj
10cHXrE+MWbrzA29rclYQbBFugvqmYlUh15AJ9YeSAwhiGr5vhHXbCgmtXWy/8H1HkaHTv1X55cB
BEP2N3K7IQzMXVd91I5A1/R4or2F9xLARaIdEm5ws4hf9tdO5flOv6n6fVipV4zTN6CMF7pLGJg/
us/1PWT6dIeQVJLWxQrPuuzLQKFoCSOWZJW12nNn8OqBq2BPCWdjYVG+v1FnQjVv55oHaBcjhDu3
eZm1r3XRTI1nII6RxnJXv8L7noOoZ/G2c+B9I+Tu4145ukK+2BGGqK5o9+tPg6MEBMMyVg4K0fuk
Z8m/trZOD4MbxsFBOvo3du3P9Fn0JRHZXD6SJ/uC+wyvl/Rq9ofklikExvf0/Jqfg4EiHlypYxXf
BwgmtW/c3gyLdx19dAZQQ/lfymkMhlAOeGvo64TBPGg+x44bcpasUmgG52UYe4d0cIu8n3UnYENp
C9ANaXam1xB41mA0vZFXEmCeveCopq/O1l+l7ATwkPutdLKmyiRYZH0a0fNfUq3PiWeHfq2pR/Ix
pYFU1SJUGDHQtGEmwjezEda17LEQfj//LMx58h9k5DgwnA4W/nRQR7my7TGWriHxRqY6w3ZM9ucY
QL9Y4hrTvh6tufAbSTFRVvoJwLsO8d2FXYrYaPIlO3gafPD3sKlvQBi5jNGuVz5x7RVPH0B/afwN
LYEBZRFwa0NmCa8gIw6Sc0Hty+Xg6HXdmQUJ2fShOmiY5RhXeEzTQXjorNNup9zE9KYVeg5Ahuf1
UegDz8K/wqljAGGWMKWAi+ZcR4iqb6NNrv3kjzYL9qcBRNOIIpPASluqEpOL/ytMu/VdUPA/WxDm
osWZXrZHY/2Kiiw3xfkTrWGY2oUaM9ySjxLs/MuwlYMomcw/HrKJRGGPveE7uVxlo+cmqttUhnZ4
fM7yy+U30EF0JhxZSfCEI5P4i3COYU4PHJQeLAu7Ns1ee/EOywf2XqpnpJ3ity6nLyN0wNIMGp8Q
SNSmcsx3NrxtcNAxO+XepeQCQWEZrRaRpuTUKmF0TV4X6oIOktl/oJqBsHRS/vQOV2CzoaxUxwPZ
9CuClskf+GdK+efqelVbd9lj+y6euzpuO2h7mCLG6XEQPzgpmSfqwQ/zlg3IyyH7z+0AFsF+mXpV
FkLIDbduvUUIL9NRwOw079hfu9M/nX3ulOtCza9KwUUKMv4HkhFEvgUC7nXgcHX5CBfCZjke/qoF
WMAiqSsoZyOvigrgiOmyL3bkNx97yXbGfitRNjyamzS8W5hD8BJ7QR34FhoxlxPI8plaFyf+aqCx
NdibMBcgy8bZ5g+zPZlodMY9+EmSGVEuTYCgNl7YnkB50R0gXjXOnP1UQrCH8DeGjOrFMLIXy5l9
XEze7HIvfvJsxMXCB6WZF6iucXYiFxrF+LV9OaEWXLwDHTgfbwn5Cnye1IXdzoyCVXFCap/KHVwQ
M5eH/CCiwxF9AzKAZi5sbBe3eJkGCgRcSkYwWSr8kww/oOWzZ/FN6vvau7kCirlfb/4TqgoAQ914
hInI+3KrKqj/DS87kB4khIC2pm1q9bpjwslpIllMpqVR7+OvG7PwlQqhBFUlwJynbFK5rZdMKskM
4j7zyfpveMd1RJLp9NEuADQtt8OlXhh1MBSGtRPJ/vUqCNrzxCOoDkC9pCFYKTCyQA8o1H1x8Kfk
au7vAmS1jOWpwrWMhFzAKbSIDNnWCHfxRE4WYz8ihOwd6m4Lns7SeDcy+otnpw1SiSNHOxHFepuo
b1zjtp8+hmeIsUcLtiZFbSVDvPXnG4pEmAp9tguWUMh+8J4wCY+I2xfWwI4bRMA4fpMpF7WO1/Fv
dHmj6z13IfmbRHrR0Za2QYQaVtmGtvlVntehRZs4xj+hyBNBpDGbiIaM8ttMExPoqpUFN+MKrwds
9Nh8QfOnimtCt+sLlYXYKasl1JY4PvQjwDIx/QhJLijIBXu6jNNoGxuegjlS/5nXqIrm2keji5k4
nI6o7mPN11FDil9RougtSHXw6QjhYkcb+MVHpvLWBVjk+0dSLD084ANReDFjJceCzCwRvpJSNTep
4LZcouBLUmXqmU9RrIrCgub5kFQ5yjdWC6dxxYaxAwzC1ZNIHvSSR64ODtgn3OHwBT4UDKBBbXJo
g28E9acdOyILMnNg8sjWKmQHFHJ4Rf2F7noZhyiwZ/0ap8SRwl94q3MJsxfj7cKq3Qx2gFQpOX7V
T5NGoEa3Q+C1jb8ih1swMz6vam+Bsvlz1ltRHFK0i/duyVtBOBuSDL0DpCdRIPtaSllIub9oL4Zz
SwAOEW4IVUyaAjrcccnpGA4s5k6dI7NQ+Tp9918F8D1rHbz5sqtI5w7+wy20sWSaK75eVBkZGuiF
RNgXQRNPfZXt8AgZm6bAoolh+K1g2JvanBKwyKCDEntMTjOb1SM7jTUKtjd7FR0ArX+tqXtjOPiT
GS9JxbFF9xYNMbXoD+2X8Odaucd6ow7GgRVAQ++vrmuygYu7bdUjOT8hrcjadsBba12Ph3oVCUXX
AnAcsKa/2zPMphZIgUIHLhsXFVB2RV8OMedVMeMRLCXXdD9LNjYdHD6f2XYOwMMJh2vDbYETSSzS
cvBR6VDb96/h/KV6eG2FwBYtlEad6qLzlczxXpBS3Z1Uni3+UtSIT+A03RmD96KAJ1sXZPcqq2Vw
xSve0Pm2w+cChoLML4gmWNvqZ+XPRK+YBpRoreib5nyPBIJ7bnQRPOHsjuM3BabFAqHFXOQ5oy1R
aRhf0V4uRFu49S+9zpGbBT50iySwyATEhqbkRN7uqy0Ou98f5RYDZaedyDmuDM1ozx5lWAU1pyio
HvmXUxPAckSbzBstde3zfcfGWSviDHGvBfKcsW7KmtWplkpyTmqPH6KzkUJiYUwjkvsjPtZKRsDb
N5YBzurVF9IReC8OomaJgxyD1bgGRRtfe3bu4LQfkM/M1ieZ2Ad9BoOsVz9j9BADiqxGkfHjRcd6
5RccuuelbGRaJl6mfgfFSB6DPX7ouo6wjpLEh/bS3CAOeCpFgjgYR4O85Uer3EbzNOTcvbBQ3sjm
mFrEF3wvTL1PJnhR2U9kMhURVUoyHIpoT23Wnk0HPusYk479Fm6KnYNOO/xgQu7Wkib0yMm3ZF2w
hsir+rv1ODIZsuqgFPdEsQM9WRiOo4rWEfNNn0OhBxCl03MexPS363PY76keAJHSRWPIfZi/IdVs
+3Lb6/tcsJ8801nel07qkXFHX8Ymhhm1LZlmzwbL1E0WhzSJwv9V/H7uBDFp2pyW52gjm0SOWQmH
QoH02DOxmJfs9FpfWszSCK4M/arBCwd3c9YJs833gT2nv9QegAhmU3v9D4jop5687VH0n6bagHIr
zA40m4YZf1rr37NC3gagT5FXmOMDFbdw0HihyzRbrCu/4vwh5jMN8zKbdm+HYG5pQfxDEIMC6JTn
4GzHktxOR911dFdawYKIqHSVI0tujIb/HMWAAyh2w0Kw9KELzNnESwJiwZ1pT1LsfaM/DmgcNC1P
EhpK7Djp5p5HdIvzKrCizYYqguDfUDRUlUZuqDsxHn9eKgvQcO4y5F58Gbw/Mcbc0PtDRznSXhDc
lqR29/DvWaOZPsRJEl/2c5Mnm0YnMtu5aaa85sBxLvGaDKxcyoUVxWI+5+48eyaoUQlr0DMZk3YE
ps1YMGkzDCfJWzf5rJJ5K14eUwn0h/Q+nkuDIc8JBrom6wE1ssX0Gzuoh8p+JOQmBW2kU/ngoLVk
9oF8Nc0LornCR1PaXzX1ZwcbSyTlOsyzkb6E4aPmXcdw7MI6iLIUPE5HgyCEdqPeMfIvpe6F2+fS
6fq0IsbZGOv9xl9DOhjx1i65hXdvr2YcW5NgGJvcXyVe2cLLhoZfXGQCAaUUkR6n/WDcaq1M/o9e
fQuyPZqwbJ6QBnuRXpF2lJeuK6eRrH5Fdd7kMC4s++E0Eq4zhIocPgX7gNfLG5WzLymM8C9Kd9lI
cG1L6KVPPb4y6cKCpqFZILr+m31FnAGcM4VzMEAilJYjmpMWdru4KcQ+Beyv1+qN6rae6v0Asob1
teLBvj7/i0pqopn+G6DhKJ5RVO1TmyioUFGb7Hwsv+zfGvHML7aNfhJEPDyRPy7HlziXc/+VwIZB
ogAZn9Ab6M21XsF79UsEKkYQceSPvsIdwGfmaurK5Y4eEqHvQBnYxYwkUXx7/2c+Qt9GxD7XHqD/
W/ZbaIGMWZ1LVC/vqcCtBAaNGj+aoGKfkpCC/rPKT3vhJ8BYmhT6m2nQa3beMonfbszibNWOWh6x
LZRJ7xIq5xU1jnY06Onabit4AGVROL1IWGes4ZyWTZvzIpkwcPSKN2u2N079w9cVc59wiKBZFl3y
luctX7vmhsiJ06bCei+ywJSOxoM1vvBoNMAJgafam0kOTfWrHajnCCMTCSk32HWtJJjnkNg8gVec
lS2jsxdWXw0qpPgjaDgnvfiocRkkWNYFyLacUQitHI9X5vCowllw7EfwNjiKjD7A/Tqy8hf1A1VG
z7iiarpkHA+GNXpB18U3bk5j/MTANFoBGDjC9/M3nZurTMH4Y/BcDRSUkNrWSERpzdIXS5uG5/Rv
H67gJFYWKuC6AxcZhdnAb8SL0RHtwaUhayg7edCGVXdqP7A/wQHUq3Ve64MMVi+MlVvo/0Vr3PFv
C4lnvH9EGi83Wd87XQJXtc6Kr9jpLGjfBlFHsjC59FJKx8xnZqod0MjcBbFfudlqkbQW/oZwNl3L
RFx2U8hYCvIcJ6gJ2/c0QD0NcMDpU5Bjd1Yibc0/ZfTHH9zEEhMEyGvGqnOapE3itqZdhAAvSU/t
ZEXp3bgs23Vyn1sP1JMLZMwDJQ3vHKEPsVYIuhXXA2rrhC9nn9BgWfw6pBOyHGvGl09m86LVdRlF
xVEk2laEn4vmbDqXgSE0wI7X3VQNcp5T5kLtoP/QR8ZUDayp6xXYa/wWyQ/RpmJDleycCz/gGWLF
OYSww6vGXTL8GtOnohW6K0pvntP+Y0VZC3yHX0l5ooAGCbj3jjdiHxqVRZtJqVwSoci0lHYosIaY
kxH14a5L32HNh9oY69puD6ZPrhVma0RqpCCUbM80TQodTcFp5kvK92HTVB34W+rM5G2dtWt49zKz
b9lJmQ58RgPNXLKOtnktkdS0ZgRfuuyhbDTliDOvZBWR9YWdDX52OvA/Pecn3MSAe4E8QtgNQK4a
LNDJntqC7TT7YPh/+taUKrKdX9VzL+8NWLbrGcyZUXpPdkXULUwdOkZZvNj6FDyCWx1gmT2VPzh4
UlRgx/JOAALmUsHGX9SlsbtVi6iVAAMFQB9wJNMlb1sVn4dIEJC6yV4lrtysM35cQHxu2xM8Mli/
0Nzpy3TOOhi3rYFW5zV2f55gyaZKm4xpgnQH+FKmaGLFQuDAV72/XfgUciUw/jloPY7tju3fIhw1
u2y62zihgM+TqWXSBWUv3XMHBu35+lVQ7P/MYpBOPh7CjKmHqB0Ivzr56+VUp4amFeXtqJf5w6oA
rQzfQJIdBQNJ9CfZuFzXz95MLgJ/a7Sq+P9HQoTvCfq0q7rtR2tlujVN96qCpemLjV9ihcepqZed
AEgFdHUD8seT1ZW3U2HpWRIk24l3tWaYqiZFXDo6WmXT3YzfjVemUqpbX6H6+rBHL8sE4T6BswlC
zK+Z0woFb57PWP9avQ/gTvkq+urbrDHn2KvvjroJi4XGEPFvMNyaULKvAzrNxnzzOr/unSdaNHUa
2jiQzLTQHfziQMFtmIqzDNggr9TWe5wkdD3hWDZfdnLPwprP9+wV25sZHawytbQRGl4WlMOteAK4
h9fSG3ZsML42f44lhLBZRiJbhlqyu2oFNDU10zcIHQpXn0P7jtoqmK6o0aQZiy3775KmDcOhdHla
e2zdyO4HRPLl3AGT7tTbxfQ8yi16bxfJ5nnkNFTJTl/G0mIqG2a0L9DdVVPaOLPJyodzCDp03Z6z
H/lo64eV9qU1oWAw64lwQQGKXivpWaQOQGZcx8cxS6pVF9gBKsxvYYXrJIVewTAFAOcConNwabng
7dbfi4apfw7s/qpPKat18ouEzZkL1Xa0lbPWcZ97+FXRKB19Bvcbxov7b4p+fiYoosS9nJqGpGqu
+p0oCuecG+z8BlhAoxgZZUnUK8Cvq/SaUppCbW9usiUD+Wb2kv4l1DaHLrr1Po9XoOatm2nRaySA
OWcIg4VjM3ktw6038Mgc6ph8IUeJAU3sDvvahHlu8XBI0qpRI2BUyxr/aS/ydbokQIKoTuKO9uXD
PWgwqfcioNKwVscL1HvzXhbOVrRaIdSzmWXeCvcyNvdNMbahQR7o4FbEyKWXAHP7zqE5KLGDm0wR
bscfJYLDLH5Y9q7ohSWV1XwKq9AizcAy2q1wnIfFoowkbG8ONvnxFDqxefncgxxF66YjAOuKGhxd
ulNFzFBSt4TpgntiPQJYE+yx1TVxhtkuGAPSwSUuBytngOujvJAIbsXKpvTlfcG+nD/7Kp6nyumN
kT/bw0GYQgt9ZzCjNGhO87HLaUCt0zK5qWD8MrKANzCIDWkNspRIjZVx0YdcsIvzJb34B3ezNXYp
ZUAHX2E9G+bquTlwcfoecmT9PHqRB6pOcEU59Hb+a0p8OpssIfVRHPD5j7PnWbpKdLh5nLAyCW+D
leImgqjrkW68WmIt1QvjmU0yp100R5L1fuVcE5OovwCOYdRFVigm5zwgx0onA+cY+xJOrCSVeg0r
39WrC+rjuaII4wUVDG6i1elUG9UXFM9ersgkYJ460Q9323Cz3UkhfpKZ+A90Qv/Ry7afJhx+lw3l
CD7HHPoogFPsII7k3/bMwY8YEGEho3fykJ91t2wsatvikFTerzKGChdT4XjhYuu0Wuh2vLioMmcC
iyO6UQKj6pnintRq4L5rcNmuyFiXSMRpghxphyDarfstWMRF8TCp31hCt7JQBdt1r9QqtgKWb4e3
Fqyc7ymo73BH+a6E50tWvjuYuH7SvcZDSPLPIHUfKpVZxqBKBymlb2ne1HuY9/jaxj6B2Hu1vGk9
eiWhjMEycxiavj8yCg8bu5XiJErqdkVzwiF38ly/3Q3HTImYoFzUXXCCGGqfqVBLQbCoYqXGBLZU
zhL814COAMXt+DaUwzeJGHZeoT1EYDyrMwrE5DoRF3wSLpGpVaDBi7knxostrKbge/mmp392knEc
3YDop6+QP3VfbMgoCccF50MU4PXJKZDB+UDjDc4cKph7Wt8KTeeKBRwoPqSOMJD6jVkrpH5Cfuh1
8eRcaJBrQxuj/ect/J2VI97pGzW7rysnMgnaCTuKYGo6UWNXyTYeXkCF/79VFQETi7RTlGNnQeEz
67RasqKppJ2o/kqvKmnhfvKUmEQOLlhrevrEj+w3/ITrbRyLx3piOHfFajGsSMKlwJPYHM+L1Tum
6lWvbAVQX26OTNUWNIefZTtF3xSE18ob10TzqaISg/wNNGId2e5LVtPu5dvElPJ823VfD99exgHX
FUvvwXssX2tGQ3FR7J1YPEwJIZlQSGci2y3Wt3TCuSFI0f0kDb8ElMDWEFZv+M4Y7Qzk8SwetJSm
8JBeFj42yybfijOIpypCR3hWLWMyD9dGQsi9t+Qxa5racRZTBKuRbktPNDisppt6Fi8oXcUG6pCs
YG43T6ErFNKwAKuMqbP4kcL/lZubZIaznv1BoPytd161h9kDfi5uI5s8uEWJ4ZUN3tY/sHOG5p4S
6kboC+un1wSu6ENYWYU7VpLGXuMXIbF5bZmxcjUPsMtegbwTD2VU3qPpXUqUuIk160XiPetpQ1p4
0x09Yg967w968nMi+yXJ97AX91K8Uy3gZKdZIn4LI62+JJPb2QfLRNn/3NuZTJaw1FYTqq1p+/6e
hq0i+iO5xaUQN4IioMuePD/EsEe9cca5dfgRbmWCR0LCZ8tCuZrtrQ90uYyv7DBKwY9OKezpvYCT
0ebgmXmPb3spZ45hYuZBEtkg3o2a73Dj1Vs31mgRhpJvp6bZnvlnuZ4p/tbytIMHXYrot5wNWZVK
MOFv/sp3EFAW7jVfqalzrXS3Ggeh7IAARBZnXtzS90+lPuBzCHpJL3b6Wl2XVHMg/aEOiThkWI4l
QvuD8zrM+eW8XVuxVsocvhGqonF4d75jh6AL1rUYxgIOdFINzZyJF2moSPlX/zmn+U3pC+NkdLPB
u/JSYXHd9DvRJFo29v977IRq2yIvyoWpJ7YgfarWiZOoq3Hsl9z4a76ousBuNYTAzfGr7iY1iNj2
8iKZPu0WdP8wl/YqiW1I9VraP0GrNizGOVyOAp7tGWkm2UqH18pPT356VsRSBc+EGeRwtkDxp6oG
FPGmCFVOZ7NbRWrm3EpDj8qSSkFqlth5WvYze5UBaeUrK6B347lpFfRR8aJIrEkvVjmX+qBYWWja
gk0lGmTJY+1ApVjEO19fRNMSyrhuuLf/NhW6p9ZG9KhqYtvZ2z+ZeaAUNWxQgU/q6akSlheSj4a0
e9SNe5WU4DvJk6B5+5sBUIIpTVU3FZXOrTJHQxoWu3z8BGMbfaiwh3yWNutLyIx5SMh9CfQIcosE
o2lu7qLmspl2Far48zqyddV6/AVDUwUnJf3tRGgo5LPNO3So/x50toAayb6OG36AypZpStCFxq2A
IADOstX1FrnNNT+d8BMlRbtOIARsGA2kMcD6LDuuPjj7XIIChgTeO1B0dNVzhKgBKJ1UGmKXyu2W
UXB+ojYPEQlzS1M5j5rRZ12hmQ2faEFWECX409uUxhxmIwXSHEBLr4Fice3qZgERTkjpOdQVvxsl
Q72IEQTqoY4AS6dJS17TfgBy6wE4OZqHd+WDb9cdfq89HlsO1Og7zDGD0lV+HllqdjgzuM4oyDtd
u+RNrrLWehFityAUa8dX812B0BAJFQ6m334xWCMw0kUJ3qyqmWkvJVvneehdwiYl2j5GdpRGW0xu
ZReALCwNAqsUqZQ86LRSRdGUxGTdJ902GTc+fvohcX69CErEs1ZmgIyW7ku7rbqibBY3ZSx5CmMO
EVnbXCkbnja/OIr160KTO3OKdOtlRFY2vzFI94vDaWw2g0UcztU+thjmgT6N0CUBQMGiU+QpTGGE
Cn34Zob3TwEW+RDX/2JY34fMnbvxwGJQw1+Gh207eE/tgLZDrop0mZuep7dSnj1MZIGlOs+zfn1l
/iehHurya2hJNs8UbpXHL+iCl2SIvRSCNHaOQsjlluHJ5YyTZUj3G5XeNJshseO+qKwJ3FGNHeZe
jXmz5pOkxHR7yi5MDnyebddLKrDL9wFhEkn1DGiint/wOPWhBzgUAKbwlV9fJUhWFzyP+8kdYBJi
ABiN/hyX0kXFG03c/BgpVjTBs1T77LglY86/Z//OR1I50EI17MjUjKxcDeK7aTdV1poPKgifTnCn
MrErXUbYysWG9JsyCurilT81h9pa/DYo4S+dxT8JscnzMD+nJ2fg6Xleb/dXNHhwqhcpzcL0cfJz
pNciUaQm3Jlv7HbODt6ERwKthA+IXAxKZyDP8qcTEG9QSLtc2DqLGBezFN47ndXn1jA8cpLC2g/I
nbk+wChPEFDKMTDU6B1kJDlN/c9zZDCCc+IJYXAuozOzfrDm1yLi5nFAgys90ZQWigGkSnhSUeKH
WCref6D8f1fkWz9Wx6zmvYL2mpyc0bx1B50A2b+1Hi9wTGU9oQxjgJxVHj1uUDSlvTJbuX2ETv1T
tNaTtQ/pMtag47H/uc93bTKjK9/AqMzMc96mSdsJROl6oi84QgJDCLyiDgc8KvjwdulZ8Qeuhhnj
/2uL2JrOXE4KoeNIvAosbgEyE4PYpdWucX4D7UYBDbZ5mBwNrLZlTEgL04IPf/0/xoj0qi2ZjecC
Pf8LcB4WEQuC4dQ5HkjlAkmXHhbKhqQaB7Cq4bXWnK1GMmx/slBUZq/aSQzvj3ejr8pimtzlUzY+
zDss/XQ+c7WUr51mmm80xRGAmvLBLxyHBJwUvJtyIrRMCk9YQbGdsIAt5uxQV/bJ6cNiSLmgOk/0
y6V7NLWJzcXmJftsTXpJuvwwRf+k30S9eV0hOouAjzIApfy5hudX1532/wtByFd9hBPfD8vUHjFn
acsBQyXvD0jDqgoQOX5o1P3GH182CgUsX3lBcqMzRc5WwUtStLbHpRUPSsn2OuzXVGV44TEfgLZm
tFt9HwoLkUpoRdsnJiIeJe+LQ9rIPugSIYNsoK4bSzKqDemrk7iWb5xsf0MhAP396lKYafflGpKk
hVBkT5p5JJaBUE5uglIYrZe+/ByfGqjQ/MnqtUXpJffewYFg2FU8GVHE1SwZ3W/dDXg+OUt+k2wd
7/89Bl8qDuZ0fjOXf54stPINyFuBd9pTmu90OM/IZpyrKVuXtwPfexXHlAUPRg9MmvvaQtV2ZaRE
fLgz9ZW7GRkowMgcOupI1YTTwub0M7bIrmbpxiuRpXI9c/0kRbNcZCfD+WTHuTxy0lFlB2bDguSD
OCB0MyBxa7ZwiSTe8fwje/NdPqR5ZyjBolFlvC8C6ukvMHirMmVREKx877dtPTPNxDLrOjfa3bW9
zUcW1fPJKvEA5drrqte/CsYsYhUBeQnCHEQhwDTQk7PCgfpTY8qv4OgjQ8W5npDGfX9MdsVnI/pu
KOnCMJuBTeH3v1UoSBOtfX+L1or6GDCDaLQKyWgP1wlF2OyvWCsW+1mSa98Qjuwnsqq7QnEsjubK
Q+uuXc8rSr/TnmeNxmF+kw9rfou416pdWszsOKn9Tg0z9Lonc6/SzqhT0I92ZhZx3Og7pY3zl32r
uX4XjjHFgK9Y2rd5Ly6bDk/YWyAtQRk6irSI/3NgxMFF7SqQ96MKVzkDysvYSh0kUmlTwHAsM1KK
8/2e/oYywhptQVn1CVW3kmXbvPBZI75oyrf/1ASEFe/rcpT+AHQW0oi9TEcmO5OBYN2iV8Jz2S0A
EHVmzEPFjbkXaQoxzVSint1hV2Avkepv/tSAVfajk0RgJXsTSQVyMRW+bz3RcrLYJu8y7n9BY6Jl
hrblz29I1Lclw0nNW2Ds0cd6DXOh2vTCNhNxa/eNfWAe60mBJo/P4yGlP1sSAoYOgRJLhHtboIHs
WiD8if39AA2A03EhXM6r+jcJIyrBu5YwLvqHq6UVxEftuR0Z6WXesmOK9DuLqNGfRfyTU17v+osx
DcubilxE2tKfnBIYYnS5QIhDoPsVeyBr96EF6p7JP/SleIBIXD+Y8w+zr3X4aU2BiOBN8+SOlqpf
lH0nkpEKXP+p2err86qg18uEL//LORVVB/klu92WunNyA9Mr4ewnGLJdb5qdq4L5NtaTOedQp/pJ
eAVT/cZF9JoXcQOxGiWL9yDTp5Fotk4jK9yi+Q6m0Y9SDZ4VdMtI1pkvs65BMh415tH10zaCM85l
bjTEmYIz7+Zx6oppnuVEIz3Bw8SDuUQTXKw5UkOFFIjrrNXeh7kO7cWAqaVo+jElFdjV9IhYHtFf
31gpdB/7FMEgrb+zvbezmM+ygUiHx9W/ealt2uKp4Zh8ISGPu2Mbjo7ORHwV1Q7I0swDG/OMEur1
wpR49UsJXY4+7xqVtGUXfZCWYmWA0BhdF3+sXLPRYb7E74PeJj7NIm5BhgRpIfSk+kZJytHMq4HH
pHGjC9gpSVFPCeDUkdv0YxnOkOQ1avfLHvir26RGYoR03NcsVXb4VHACHXueGYgl+1klXNbj8iQN
HU2ZdQZATszLM3BEZWsy1AWjUsWqpT7qKd8t/dXLk0qLElSCfkOxBWq0SsFxb/zISZI9Iy4An+CX
lxpm3DCTIJcH9Xbo8dQ1NGeRzBW0CE9Was2nIbwhSuZUdWL9ihztWl1xZubSIzNP4LJsK/ihTOao
SOrOpuk5FJtzzmn3Zmk4MfcEUNN631fUS2OFDxayuU+fjsZdGOvu2pCrvxXvfVm0peilwHqFfoAI
30cfB5fQ7RjwUweMyGw04QH/r1M2ebmyuU1IKQgOOf6tUXkuM3VBTOGnWiqxelzOxlRhIXplkNWR
l6aD2tDt6MvPmjXGXGCcQckqL2jFJ+gySJtFhOfj963tMobgt53LCLLMMToSpxzscQds4M1ch0Ww
lFtdN0jlDKGbr3YOjRz04qJIX597n4/rqGOmIjizD6zI8uMNutKDIVbYmOnZ7KgUhBPcsRuEWKlI
7ACOHfa6HCj3roI4zm1P7Sj1eAylGtXHUTNXVpprnEY6RNnz7IA/r61ktxnzME+h1bas61QV94qF
Ufd0VghlAJvrVSc6vFmLlPboESeO70tSX/01vH1WFW6YCtDdeSoPDhsHGVqoAhMTiLx0XHB+eVQT
8RqJ5+VRT9WwU0n9C+AmuInELKXlRxdsKGXUcyIqBqZ0R4DQnTQDvdvP7AhorML9N4U6DT6qBMvK
0yqrZKd1mVtIxhrAI5VD177VR2ABrLHTDpGewgRwQNgUpvIqvyI3HD6wftmSfEjBqQ77d6YvcoSu
wTwySXveAWSzrxLmvPzxc+Urm6isvOTZhqb3doE8MgZg6aUU/+ViNVOOvioBYG3+q9LRUf6NYDQw
d4ajb6YWQAxqcbBcBMLdP9yhjWQT2vqiKILArpZvyxOGVLmmqbogCFsCy6ppBCgJsrSpZxdFkJcW
hkKmJy2qnxbkArydARLUa6QftzvUyWZ+ATdG8o5IvWZwcHuuxB+5FMQQi71RqqzoLABv/F7dwAPN
/YTzdgDN8X1LAvNRbzDCvG8tMXtLWAKCgJAODWTIroJkpknZFnZ6EoeVDUTqw/lV1Yt8e6U4lkM8
LarBUzbS21jBeHDs9015OKoIaQ4IecvfrdfnQP+IBWAAzdnrGWrmfZDAc3p3BAXmsQS33vGMlmTu
R/FqG09bkvgOgStPoT52OTe84nqUZnsGxfUHa58/QoSLunDZlzGbve9Ysuv1szp0TUsrWtfHhItx
adX2SCHRdO4R2YoIkOLw8xf7g5sJPOltzdKDKrF27SkPSnRPNsChe0zmql0RB6N14Gfs5cIOykzV
itaGtPWXYuO1HNId4E90J28/7Es7PDNOKuSIftiqxQPxC+3YTIYe3MWRT+NDc+f7SR/8TYMj4n3W
lHBwDOc0udkyP1ur/ApIckXFAv9QuTOYb49I6ZFxwGU/DU/PYWPVcwOCiHIbPeyaLyCG/KFPXJBa
y/7lg+QC63i5bpfcbKtQcd0V6guMTl5KFy4GAFl17G+GCfIQZa8WTT0QbpBbb0ooPsottLpi6nzX
LsvJG7Z07mh55i759tpNETisgULzxkvQgNXsb2FsUVEY7zV1lSYipJNbpl9Ufa4glQzx4prsahv8
MXagnR7Cxm8ZPF1WqDnc58CAW9yE33USR/GHiOGngVCAQkA6NdnuH+P6Na55ML/Bwt7tlZkVmCo6
s4JMiQ3HyGNJOzdLlHGEJj3amclE1Rj6DR2/a0HdnmQgo5u2+dR+R9o4Kq3kCcM990XDE3bYmYgC
TWUBXkXjSFBqPy5msPxywcY1O3voUdwlGAfV7Q7PZwbsAf3NMG1FCKGRMfGX/Us6uD/PnbUcz0EZ
T7UQuDMF0QQyqhI+NGBPGJOSV2w80vQqP4nocr3zXA0SmGal0kGi6KzIRYWO2Qb9wu1nauoC6e9K
PIGpU1RzAvXF5TTqeofPWbyOnXpOvriCHA7sY+2156z6y14gAlmijVIjnKCZsMuzd5YatLCY5FVi
qDBSFwWwfVqEp7sOHm6CsX9MTJdAHOLsoAwrGfrYzHnI64Z+dGPBdnnYKpkZ7Di8HNFUp6INsvjq
bdIGEeHNo6shr8PcMBRsVfhLqJq0564TJfiNE0Qtz5vBNKxrORZ8zWBzV/a3erkXKZCgvBng0YjT
ahTG1btuJuk+lFTAY4UJ2TK34i/7WmF4bBLj9VaakMYRTGyLCqId6cPL1XspgIpSsrAIIRJeSeIf
UUspwUsK0JYbk8LzKhzHl4IXbFD5HAvl3JgaxYFMWZF6Ju34n9zMetxzGiXIzJxbxakktcEbDvLs
CcGOL4RivPLDvYRyKN51re6wehYt56mcMW7mo0azbkqb18qzO+qNFh2ryjQpzQWB9CiZTgkPH83+
xIGqdayRKoboq/wnsGbfyMLis4bgAFQazqVC6//00OH7bCjVtJcpNYddH6yt6VPk9hae+LHRPOyN
Yc+EBPaggO6tLouNgO63JpOXp+OhV1k6AniFEnU5OntuU+1nBmAHtpu1LVI0ofX8bwnkrYHZPG+m
Vm584es2tqQ4WCtPMf64mcTRZtQEs1Ru1fUFspFQmXa/sjb2F1MAZDnoDxPtNqz8wSzE++AO+Vv2
z+vEScgJs7rOki1CsJG0XZc12b3nbaFlyqslZ+qLorxQclRyZtsklTehwy4TzYNIN7x3aiGRWhht
wCS9XIqarrewC5q8s2PxY/KDV3eCjI9Z96kHgOtWDhfVsH0Jk7u0HldpRKzmOJN5tGVD6V986kS2
ER7zSqkLyLTqdfRKbuvoaZKJA5RItDuBViY/NMoeChLndVxyGlTKMUI1FdZwwmnTxjwyPetnhL05
SYvcGyM5PUi2nWs4rELG8lwQDf9cQX9AuY7zyM36/NuFJUs4wh8wippTkrCAYR/7uiL7inO4MbRV
PKA26PbPGuj6SXX2cuH2ks9tYbrYrylqMwdg+ZPe/XNpq6hn0ynSsfGWtvvnu8pKwbW3dUEZQvhl
s0LylDZavxgG+OcDZqAkZ1ps43ATfOFUbd8LS+xjQOrZl53hOittEMwHqnsXZVPGYnZT6re/hXXa
gKkfuPLvQAee+Z+/yndDfmfNuhUfMAxTYpoVmquP4zh8sj2vAl89f4T1TtYlyOgQjAutP/PCdxx3
maMdkYCT1IVyM0o4O5rRQGyDApVsj0ssYtjE3PUsuGMCdr9ncpKbso8hOx0gWJP8zFAHtZWT32W+
EulB4c5qXG2Rhj8rcI8UsQ6RH9vI0eczG/5oElHnmQghD7jAH1DSjgGyGY9KAiLUWvQeuvB7LoXW
XC/h0oj2JOHux8mSFnb3+wdT+SadOEpdy4hiBvXyvo6ltOWpI6TncLUTI6zhAca/BpVBPGSDqsAn
3j7E2xlNsBRBjSSIIEfYG3y4OnoB/2R4LHtb3GOFOBTm+2dD5icW+blhm5O+I4Y1YE1u/lzfPtei
FX0Ie6Igzs6do7rDdFw+naON8iXX9Bh7nLPiICLcbqmgti4tuZxwguk8PQ/2nfSzrwNdukq9HdsP
esXaiiT35IdFpfS5xciKlcxMYX/rc/u89d3S482jEfluSan+ziYrOrpe5g1G3ECZ6csbIm22etKW
QqULbw6q25rGW8SUxR0vgAFI4CwRiLtGe1/Ie5SphqkvUNvg/w0BOfVylBBTcvZdjrg7bHewrcE1
B2yHneStmkFmZ8tfb79iw4reLHOYv5qmbe/fgHJocgOkzbY1pEr90Tn0Zt9oNDXEhu/KABH4zwEj
f1Xwe5pRr8StG2gjMe3dypESR5K8sE/ulvKMKVofu7hs2SNEUGX3NhgsE2PdvU2zWO+1Lgsttu7s
DhE4OA8P0f6ZUybV5k7HcDq518q0r0KwpGrC/gSqB2dW3KXwxYWIZ+TaiUOzHeRv6b3612hCoONH
CE340JMM24ajW/WrLjTtHg0qrwjcTRe88LXDJA7a3lmylj11Y6eknGJAQFmhpUxDZxVgdw1s3WQM
iI3PSWXUmXpw8VSB+YX6wJlXlQBqfVyNIG/Tl48iFXRyWdNYwxj5hsvrIiffQoM8TpuSGDfitQve
TadRlfKR/JaXvA/z74/Xy3f2jHFXo613HBSKibNVRaQY6YDReiFAsT4HENP91T2Qs6aD6eZMkbwv
emX74m+OpszJrBmFrl1OPVZSasfXpF/pLtdQ3oRA9ifRDU6zuxDHj1SDJhLrpn0ZYIqdF0ez21vN
qjjBjruJ+70M/E2p198z/lVzpQ+ev9QOj/c2RWLLRRTHAN5NyPVWDFUUTJOQCLha+XxDcKem1X7d
yUyXfSslu0E7zsMv6QcauTxd77goqUohDori83/GMkCQ+8/iq+waYB/dpbT6XQXXFeHHDOPAuRKT
cD4oTJwDP9uCLRinZqJ4mdOhppsS0pvsgCGqrpnQs7BhIr9T8y4//NaWSMvOLgymYbJnE6WOfH+s
VqJa2/J5xRJFpb2YjHnAAdLLMrgoxyfzLQ9DVRZ6Ut4D0Ijs+8zTdPdQqa4fD2FHIdwQOOM+gK2J
MY+Mw+Wk/n6dyMidyqlemzscDD90YQOEludYb56ZGIromDwZsS2vwXtLCK+MMlTA38W/VXx/U7iK
JD78lrW8z2XXkp/azM+D2cOU/Bc7kmeyIRRKOP7J8L7R6KczZiUT3JM+Ei2W9R8/AFROWt7Yitp8
Vbdmf7ZsKiOHGD0rBtj2qp1lTphvwssdzGhg1w3+xuXKhresHSrJHa/H6nVJylcKodYK0+ELIPL9
GoIAe3M7ammE26Bal9P16ugKOtFI2jQRSHcj0NsODLUOOORvt1V3DSc6/jwD/uEGL9am017LFRrp
BAxXPLSkA7l9wfWZ0vNOGSiQX4iFKTD6YMKl3KrfWKIEmCdd6sTEyZBHQ92qJ8PICc/4hhk29Btu
SUrrdxb9PsPmdnb7GMLLLXH2190st+UN4FD64gFdS0Mr6j2TD04o1yh1jghn4COfiaHe5VntQTvw
+/D2SmIsJZ7LqB5c6h8mLIqmmw1wmD+Bq5MwmMwBasHURljbTKTAv/wqMWxZGKxiNhZY+Xc9e5CT
+tRcgNlEVBsF6L8CrB+hLvMgK+7YhLJYz1mQyVx+1AZoYXpC2c/SWJzSnBCaHQPNL6OQP+gMRYRj
VAxba4pXR/sGt+HloVJuskZT4SwSEFUHwJPVQ/tdcpcS8lLdWQcBRgQfAFr1oWP+D748bNOdSYCj
b3pzMocHVJ68h5JH9nTQOScIdgou7bkAnPJtNzSA/VU0O/SDszHcQtAxKOXSnP/pzzoDtanZOevI
nwPhaVIxkjpD+yrfl6NLfZja1k9ya+tPePQB3CPBFjTiIiiUM5gqzpyvkqvSmH5mvUd/OD49P7gf
VKZvJv9gHL+ERPYqLuh7bLAs4VxDmfGmwoG0BryjymyljBjZn0LfGHNZyfwNzE2JxX46eWOHVocf
p80BxwcLTE2H3TplGPmE8noSLBaerWC9Kd0ugEdIK9Mb9ugNFC3+W+4THRpeN12rJxoCJ7MZzODM
7ZRp0gnJr6RQykgzD3vwvNB4277m58v7Oo3Z+6UeeNGVnzb8PqXoSI7H3KkVyGCCq8YN2Rv+gEjX
4i/4pn5mXxsCPKZDNDA+1+0gnsbbeAtM7gBS9tYY6VOpTm77OWIfnDo9dGpCztWwt/9IRd7hxjnk
loAvEIVMaUpe4mtM9YruLwuxGjoX9gC6iXIbNQstccYrBgvg3iJ5XSOlNI3XFHvBPLRn4XFJ+njW
9SNOkj7FGXuq2YpGajp1GzrNu92K7kk8x8WXo/Pw2fPTiOOTw8tox65lC/H6JpPT7fYFjTIkXn9P
rHNBzlyut2DJJyhZhRZwYonNez0yG1ujwMfTNgasgJUteOyLUrAkYaCxfjzg7iVVcbjmruKnVXqg
hW71MJvN0rFnIhKhZv8dX0ycX+7KyNQ8Xzey0MXszrBEbIZl1/xMBtsTtTB8jjWkDgU3aWJixVlL
FKKKOUuGPPqeRDKTVMqSZpkM5lt527V5hvPQ0kQ5SPAHW3461rmbseWl0aT3CWaG2PEYl/yWiW2P
MT5VvGoWbcB8aikiqL7/P2PzosYMcsRlEJmegfT4DsU8ONnA+rPNxy4QWjC7hYstc2KqkTOVM0NM
ccWyb4D93KIPardpubMa1mBSHTxug59BYJtOF+XNhTEbNHT2gRLIEypSied+3aKvYpjgwc6vadNj
7ysrlxEvO+PsCAEkNWUjp25ZVEZUkg8gsYS8bbadaJskO8dxRV+2KYhI4D6WkmnMSFc1aOhj6jaC
kwKL9OiDcG9Tmurw+D7kZeQaJXj2Rm91wVZOQUu9hpzQsPfg4N9J+XsKXS4Lisl/CFfiQVv33HQo
7lpij0ZDONiXY3YUKq8r7EYBs8SJTQHIQ2EV/MliSBitJZqINXffhpumKoJUCSqVLL9W2ldt/YSM
/Gf3doxn2bqcOlJsbrOJy7ZKkMJb/Mmg5blBYvJEzrR3JJJgQmpNfucA81gC/ArvHRo8G9hGb6ET
GDataWZq0d0vmPtTkGZcU6A1+ppSobyjxLxxJnQtDqFsdXofW9sUXW8d6TcGclKwzjQVqZqftqfv
vyuiSV2duaw+ffaIQ3wAPIWWhsWm4mvyLMuErjlhYRuJidUX2IRpoEnXG20/ragsAnbt5AXZNM3v
QZssIcZyyURq9I6WypFExH6ZwKjtD4r6AUbe4TpIC2ag/Fcka5V+Dk6Ps9fUTgoYnnp4kEVL208o
78wps9+u+NTW8FPH5XVLIn2knBU/VKDp1OxCiu6rtXgvioVmrv4VSthWSyEbubw8Cc4D4r6QhSyf
xqmb0sjc+9c23nRA6j1PLJ13fGla/sYlI941H+QIL4g2QScV6yEN8CE4Br2OxFmMgoHe9SWEVYSn
BHC52Cpv/3jlvlgBo85rFOv4C2QWZscRxnEbEnWfdde48V7gOpLe+wac9XXi9mHeqh/ATZCaptRd
42vSzgyzDBxkYhuCgsr97p6EluHrFZhRiiSdou96rshy6cK8Om0J/sIbQEG2WB8w29jy2QUepE7i
SQJHgg41veIMr2gaozt14Z0FsAtcseHfF+XmhkXvTaxQb+4wJGvi+39ZzMtxSgt4PmRmImUxw5Iw
RUkBlQ7J6mi4IyPddQ45grx7exjnnUm+OlGjG9xhPVV9SpQ2RyGT0UfCTjWnWEANVsgx4Nnf5elZ
dwlagBB9e8nJYTyIMvRXY91VSAPJmu0ANQQo9d4Ne/In8aCvE1NZ1B7C6aYb/VuSqK9IfUlvTo7i
vmGGX5QbRD2Y/bmYctpkFobg4wn7pkrUsaAHS2Y3LK6Mz6Se6cfAzYuVq5rKiskaQ/q0gTUBM8y1
VwFE5j+dDfkGvlNQeUD2vRs+ZoQnURKZo1sFEaZQ1xY887r/RiesfmTAtPwXGp4rVy/Mm4DLru4M
rfv+ZCYIGPfwK4kgtgiUpJQvMDE2TtkDwvdPis2RBsNGg+CMm4cCi8NbN+0ucnANHGy0OqEbYq7a
36Kk5/5Bhhj7TkF4xFrI8DDfmLyfLcBDP/ia1cOq4YYU5eTUAgZgkG2WhlPwzGmpHm31iR1L88Ym
J6k1pmPi4dUDaN2RNtIxMbNHo3fvyNj2yl2WWVc9XRF4jqew5wYSosDWUfilTBw+RrAn1QXA786c
anWjHtq+z1qVVVeJDz+nPzTDW9SNlxqefWvaOzBDy9ULQDwvaqG6R62YPGZys/Ophoabi4Kjqogl
lYbSed3JNsoLY2lPfgapHb254PY5ZQq89aJ+XjrQiIFeeQjZ7mG1zQDVsRfhHzJgwkSxIoFxKJiO
qilx6wMYojm+TjnewatpKYii2x1azhv0fnmYGJGnRLFqXPKpug9A/BJun+4gi9uGm6dC5Bmk/oJi
OI9jg3RohUnOUgrchaiFBIesMzjq5Wr96eHd+MKmT3+J4RdTIkwRwBcmL9SNdNcB/4WwaIcTXdsX
abxEGarMAIKTAryyK3bvOu4XXkgT8rf6EOJKL0NSSSb4HDYJ+ZyMU0xkV3b2sXEM4tGgI4bSO/Qs
2/PHL+Mn22xJAj/AbBiUpss0nmhq2PdpbNK1Z5A67pQ/TXx0fBqE8fJQPpHSv1S01GxIG3sFutbR
gw4orglaXcUE2DlIdSc8lCMbVu1XcSN86vGS6lHr4AH/gS85pkEHDOUR0HHT7J68z/xMvrg+ZAhN
JM252QALHGMpNOT78oCUjvTaZiEjmkNpgf3EOLJ7xqL0o7iCEXkUCFFzoXI5bXQio5EWBeq+yXAX
4/qlMegVPR6NZLL24ZJV70KEtqMJQANYHg4tTwIj4lpC3Xn5Yy1Gd3TuRUP0qUeridc6nMO7wkks
yE+gM17fnlvZO8bVexUnC12fhSPKyZOp68msyJ1UhwalUmYjwv53fdToJ1jZw8v4do48Iu3S3Wnx
42BtqY234EnyEADaJrc0fY9KMteQBL5O4yDXxY/MKDDGQikk6EzXoAevQeBoWsnOh8wZpdSR0azR
JKLSdGvKZ9wooQ2iPEvCj4OEau3PQ9dYY2fkejNyZnMJeZm9ckPodKZ1CnsHMEHhz+JqMJwM/mBJ
bsb45b7+9Hnfofocz4GqOzqU9vJo17U+8dWAyH6ucN9fwyc9q7wdZ6znpQyTzlNfNRZZgvftQKe6
n061jU9MX6kCY0nWEmk3OTZFmkC/ugNmLLmGSgK3GNNcAGCENIV/4mnJ74HfHZKsAMb/idkfWYn9
Kjh4sxVC0QmZ/3yCDJSoOfNxo4aLtAemhyd3DRfRlTZ2B+jiQo5Ml/uZyh3i/lfn3myZrm8zZoR+
bncTC1oXF2p5kbDk+w6SYclEqmDkdBK14QuywaGr7uQ6Z8CYOARZbDCdnDD8sQJn0eFsI5/hmbHa
vV85JEpfKv8Q7+3B9AxgznarrlX4kXFlc8H9lJXrwWvp7mAvsCI43BUzQBV2+OVsefqy4Kub+gke
9KcIF4o+XGQ9acoZhkm9WV+mTqNKe/TjziHsqJjXx69KQTzGEpGR+mxALpDWXWtsi2/FxlcRZ4da
+2W93I8T3chQEz+Cmd6thHDHk5tsyRz/ec6neH9Hms0egqFcLtQHm0WqkjYsS7l1Lzo4wnRdKfkn
/slqxwmwuBc4/wBNvb2xU1k5DT9/2ntBXFLXvKdtdns4gPp+nvXC6+ndTB5qsgUcvJUtgD66AzrI
ZUsIJqi+oWvvVhkEpvaF6rmNw4tAgpEZSQQUeRBy+YzSVV+Sa+BIzBMDmFpuDdt6RrXYA7Dr8JJ8
+e9PB0d75NWsGh3/QBgOnIio0eM8ooyF+8kejyNhh4GGnmbR3LnQW6SVLjXAI+5nz/U+wEt2J5R6
cSkx0RmoOU44aPRLDi6WcH1Uv5zca0Lx8nbL3ouNKFLdK5ZaHCCIgkzJHa1djhlQ+8oZMptfoArS
ELiGQHtOV2ipJfoFSq5r9wM78q4LLfQVDHP2oGxzDrMCmIcLoNtxvHUXtvv0iJzMwaJi5bbk2K+Z
QqRuH8ukQA+bSS518fbTqsRZdKoEsHifo0aA5Py3jDESkT40i/UmJShbJQ7FAY1kg0ZjsoHlSY8z
f/b/sKxYInIbKbiuAosrCW2Uk2S3P1qYjDfIMON7FSbAc02V/P98rKM3w06+qjCHUWFc13W6FIC6
d0fM5D9sp28wYYl8NcNmIL0WeifM6uNjgx1DMf60mvTPw8mGfk488JtRaTfOPZVh/8F5puaUcEsm
/h2ucvULkME+QF3PIoghNo58lfVIhPlSaCdUQ4ZMPqEQa82MkLNGuRgtssfeegxC4VQuL+CqBBh7
mdugWzsVI0ZhWTertzYfW9ISef8JaBzmM34BmOTesYYRs6QurICowjpuADrwmb+hLqVtDCvlmGU4
J6qhz8cE69mdcVRnkIEh0b2ZKkjDYJQ0ZCtiiqDGycdRlFYW29caRN2f6V0v64z82vvnhYTP8QWy
Tq9trzU0LnsU1rJ7tmC9Fn6Id59qiV+oWyShYbN9Nu9rS2Fr6xrBNtxrlSBv12oBbxJFcaCVmjmX
Km6ueW0YXtaADhPx4ukZHpJenALp+242Z89/Qyp7bY8Ni1N+LS/vNE1LxYq12hgIyP6VPJk6i0lJ
G4xWkQ99K5qGE0RI8NYKd/7nY7yqeEncqboMAIin7kbDEP4idrYKe3oftz4mlwJICKTGPRQAPTfc
0dpx8uaLYp9vQeapJA96FRnK9J6FErnEuhW0Pj2X+yqztRIJWFsB1/ldALZ6j82uC9FKeqdoI3yy
ONkMvjKPYMX2misvdL5KA+XNPzWVHtPzndwuUJUvw0IrnvEzX/LcjKYOUkq/fn+rPZ58gn+j4Dle
qd9QlQak6fhplSzeYgf9tILZg1Wyq3lSDzNs6wZ3vEkdlBPRx8mKNNFvtHB66TIi3e3PvQholdJc
a9qf8894mBwl9wJAVo53HaUFP384pCFpy3jA3W/ZxgoBV3w2PTyHShxRIiltJ66ID3mjzTGlIfLs
aO8NHLS7V5DLFNKQ/4YuQGkv6rNuzOR1FgzfsLC/Gk18tit1oWW+yJCyPAENTP2RB0N3KhcOg9ct
xzEPNbt0/wWHD4bwyBtWzSlzQEavijb8s9LKDKK3zLGHApkbXhI2yRcUaQiF0IVv2qI96h9EZiEu
1+0l8OYob6+eslN0GIrRcYY0mz/ZNVLVwlRGK5IE0TicThdlvVgccu0bgfhaEyotC/tKr4QERFFC
5RxPUXmX203ny/035Ljwp4v4G9BxVpKT7NnlCvQ/ymbXK34evjhnvkWriz7m+uaJkPCpc2kuuWnf
GY1pVzoiODhjLCPmmi2QluEBG7syDCTzSerUm0pdyk6IkV1kkAiIjy999FXK7OzZK8JOsr2qgf2c
hzuNDuiIvZICNZm9bfjgt8bKC6Ev/o07kUc9hBErfxERMErGPelE/mFAb68b4ZSAhlfaV4W1V8Bq
sM4RY0/VyUBcWu+ZJhQ7fv8ImIVdBFgeYtOtSOzVTd8pKrDlmWWltSea2zimq6FatBlEky/jiFPd
QH0beTn/MM4vsSsRqeBZe+BF/NMAzDafzUjVOJTKuQBunuFZsK/OsMUOGhWNRng3SettHOZrUq9/
4MBXfh/beadQGXlGj5VwnFJwgxNMmlH1DinEoG1Aac69Sk0cM1tGwHKabcHg67Tt3rVg0p7N9/lR
v3YbjN060HQuE/MhXEbof47Dmr8quUsmlWOCZ8jg0Sta8mp1Kyp6hdUr1cKjWTwNoAvWQnIlTCpB
DHmh16jRdMpmxf15jvpltKN9Otq+3EufNy0DB+WJIrDFPoqWsraOiqiH0bvRHc4CM8yTEv9G84Gy
cEeMDKMBn9c/tlt/eR6nb3JGcT0S2f+ZFQ5x6JQipfgs64WmsYZuUkDFRC0Tg1QVoJyB+6Zep9KT
fpE0Nao8UFJdjy+9bx4N2lVxgT1+aTemahODPitOzSd0fMZmbBQDkWrjpKcgcOO+7s9j2qmCJwhC
MNhmfkA7ByXR/gO+9kPzahuuem4VOEOxmzf1S6a3XiKm8qOGs1OdFBa+5+pYH+KvsMCnh/7V6d8s
ZSPNUhz+ETN5EBHJgoCa9Zs5iVCI5IuqNvovmgFjMPPQr9Kr4bDQzzOHY0KVyIr/buKZu08e6hUU
krWRhycJjSp4lx1/YSgCh2ILF8+b+Lqr/IPsoO3sf7njj6YBy9XUIHx7LMDN/43iT3R5iffh+DEB
K0b1hwuVh/feXVG44z8xYM9A/9AOKyjWIXQSqbNRBOASznNGrVEv365uF/V0Bgn7lfitTuJdkpR1
Y4UVmg3ciQfahkCvwssUqe3gaxYyZVNGXH+bHEKnmQQaeEVQ9EarZYAk08lg7TSAMDrBXn44Dlzt
FLip57+Pfyv2QYnXgRHqgCH8nvTTLCW200VhwS+QinrcJ4S7sfophXGmMcj4J38stvdt9ER4E0ew
DrxZwrlUBgKtwWg2PWrNw+K4A/Nwb4sNIXJc6POL5AltruoQjIvJ2ANn8agkEQtCrkVEiNc/6Br7
cRwN16nstg4MgRdOXDwxBbUgXJfzfM83XTLkr+LewDRL/LOM7m8c18jdkhFZ3m0pQeYQiyDEOa9O
DCzhe5k5D3eGYUmabi+Q2r0nRnvbu5BvHyqov0OQ2bbGPFutWr479erfeyKrdnBe5mFdUh+5mykA
ZHeebF7eq13EsaFo88aD3YLJR+jSOrLPqWCxGiaAt5ALS0OF5Xvw3xGPEI93QFaqqquW+Quw6H4v
BeLr72HUGzQikLZL5KDaGe50N/OBu8Kpm0vnf9ZdI0fqVxM+u94ouP8BCvNSW21Q7Dk3pZjMxFet
c/VRTejzpKfcN5MTfbolvPZjY92Bap63o+zu9fl/YMM9MSXhLvsAfIkK7oxCGE4fQWJbcn/6r6RH
ds1YsrZjfJB6k2VLoFmXzkIrKc3iaL/t3nuvRdITMXYT6XS4nhqNgHsm7mghWTZofy8L+ZikCdXI
bVhlq9ohhSn5oYHoQEzWyRBt0B0FDZSkrMAIMADwS6jJ7tSawFMlxY/bFoGiA4ZITKLBSJZu/Lwx
2C7knMHqRKSOSML93UHmUHVjTMQrYpndDHNsgbHP6oYtLozOmuIEjUPZ6/YddSYLF60l05R0dT2O
yWkeeL/RSnsCgTBWcfQPd1P2d+SVuRcUjzm8ItLqv3ubNmLXvX00k7xJD9q6Zlf5NXS5c0O5dhNt
9DhnMg1fCOcJUfz0OJg50pidbt0MQwfELjg9ebjVsQza7RrxxuHBBw75rf7CAYzlkVx34O2Hbnot
nk3iV1UaUC8VhuLGYLsAqIk17RIkwNz0ASsTaL01YTjZkOH4546/pL71MZrvSgl3dSXq+HrhCfx8
tUDI04VmMl7Oeo47kxstd5e/RquDapnCRS4TvJiTEBB+BWyWvolHwttl9m+FbUJWkaByr/bHoDmo
jPbv+BkWptcAg/EvRfvKSt5DuHoCR2fiK0b78YKr/FmNYghaUEvt+Sr9HxHdgqmVGZE7DmVX3iu9
OrHqLWEi9yKeSNv1lHB6h3gs6wCt92lLnoIPWa6PnfyMIbkMtC2UsxeTy1PogRVZ5Zdv3unyn5zJ
mfs9B3Y8kylov5ZrR89T+8Rq0Cck7UBTtBaCiLbXkzIWksJa7ty8Mba2t2m/YLKxJTIQPK6sDcpe
v5grmmUkrQJSCotQX8+P/40xXgDYQElvkVfQ80ZPI5ut+D5qXC3BmISJnj+wd3pS3Wx/IVE/mk5v
sVPeHsXihZoKbxdPE7rwcp+W9wF1Q2duiTANbKF5mSSlQN2WYlJ88oIUdxD1CfeUA7KAt/WJw5X4
dCa4ysDNU8dZuY+1W9NhM9VSvLNSoDrpUmZFm6oqLwHGPSC5yGb7qaM9oxcok0kmHGQsn7FeZFIm
YDy6tolHhow7lUOHL5f6DonnWVF4VoVg6z/RpuIGICSlF3AOOfTMhpGMJ8dHdpRR4w+0xmGJviiC
9F+BqCIGpg6VVj5EEUkdPGyvZp3iBWPj45i5XdXT4Tl4UVa5uZaL98tq85nP/SAzdHLl/qRAglbz
3f8DCMxHZW393Z2OZcBLdb1bOyANT47tqZiESUcI2c1ZdxO3obY8MpbAuxGR6ySosbSU8p6DVGnb
P/+g4+Zekp5uWDZqfFHfnQUW1kNA5kXKeS7AgVOaFHCDjUtENIqRzzg14jgQqf/uoh0VU1aBPSS6
MGYq9nCA4Dz5Ybqvoh27PBHcXyW+98CsRHH6MknGO4sQeqOiaiXtEJ9cBwLcSAw9m2sSrBdeeVMG
jVrACNMNmDufFgAhqg2BbPatml+CTYI3AInpsXC0dJrfRnuu5ir94oarnCy8tReqkAcA8SuIrHt5
HmmBvEsHeUgl+JezAVu5fGqLQL9b9NPsu4F6QWxef2yuD0XOHMXjhgc3SAbkVmEhCmpIp58u/x9m
a8TFR7U88QZ0LOPzkek/MvB4zO+S3uyf28ZtWYuG0z73hgMa8WuXwtGXp7/caxg34bIRP1YvCdmg
K0UEJkirvzNlKdOfp9sgeO5YhG3YsHpFckrzePiVAaSoxWg5DqA+yeyctyd/VYqoujBOGH+km0LH
rA1h7LCPh91NG5B9RDHoArOF7b6sBxAYfRJppKqq41XHGu6CoIDUD+wp2RTyaiL9wrFOsneBvton
/dFaekzpMjAb5Kp2RpjKMvBYAS7J7xPRlmISUFPN/URuPe0qZ0g43K51FOc7Hg0P782DzvJPVoB2
Fmnmk0Gj+kxV2DW0aHHKN1SZalMGaIJnP9hiUcAjDaMv97GCAF6tsodFMk3I/J0VzMMwhYndOyK2
OCG2ffCAHQ/YLWzhIZPf52/8GjU6arwWdFJgy4BH/GXMPHjU8gTqcnMULRFcIv2Nwxu41HttuEPW
RhABd2n19lfP1fhK/BMD40D3AhVJLhWH2ulzCSMofMSh0LwFkM5mymX9hs3zTpmCwBVsKOZH1wjt
I117N7SABZAVasPjCAtJTR75YrkieC5LPomtQrwOcVn4jZ27op4OPOxLoqstME0OUYJ0OF+XaIuN
sXUSyHGpqvhnKm7fOt9oB6ZwTpammKtDMpK9KM/3P74YzWluCy6wInDK9ZtQtzOPKetxvEp9rowR
RCFWRNAHZx03S9OqcRCoz3DGWlNENCXO650oIhgcr8FHuuNcm0kWutL3NzC3IiqOvnGaDlfXmQsT
DKpfPJuII5xwcaHHog+cuNBmwiOuPPzKD338LcDTfOOG0tdm0v3AOdnc9VUeYdITR4mJESFSQ5Hx
n66Gw93t0h233ee+N3n2esvmj5uaqU8S68VSL4HchCDjhTPbeCk7bitLF5gxO1KrAu69GltTrGy6
mF3Elyp+irdf+6G6k2wkH6fXdVsKe+37JEHlY9+xdiPIRKrz8e1tdYtquQRu8doS1gzcyDQ/NtB3
jWllyaJyz7mRi1h4+k9Uy4KWHfwJ22bAzTqHXdW2U51BHrnw5cBHQAucWRCvD8bKzJmdwJaFsgC2
hpeSf5W1wfepeVdw8XK/0b0iaB2FUt1Uk0btt0d+ecNkCjz13pvuzTh72As/5gxvQ19lAG6+z2ip
tr/mQ3/97ZBGkD5jxk/3H4MJeIDy/0iTRguBizfC0uahgbmpAEGKHDwCgzF0oNADNDJnwNVJdKw3
dFvwn9EcFg/nTKYoZAoXi1WE/f2r4vSHScmy3N35+0Y8gO4l1mWditCxoJFa74D1TcJNf3emfiWG
QORt35aDFGVmpGiK/6SmbRJ2zxYHFu2ZQ3t4ysuqddVwvEuilnjzsrIgKFxo6TOZOGLLQUoQUvug
tNlgm8N88IMNX4OEW0PkZVjhl3/GB3U883swZ7tQ+e3H3DQWpY4mpdZdAUZIKjH1udXgZB7JF+dd
z2vJq1ltldiz35C3qR7PUNXvQxldpf92T44Ohw2rSKm0ndc4qQLHtu/NA7yzEpdTqc1xX2NA/Se+
YGD82uLuqMnn+H7rAbNCDWQ+kZpM4/NeTYNusSrocoEYs0xNYKDGHYPnGczXxAOp/16NXMJC/ZAB
95N1t4JMOAz+QLq1Ryd2qKvBjR2Kfz7QLdtCr/M3mpL3Uy5X0/eESRlfFrmZ3ZPA9Q/8BVEFQdlD
Fh130KWZany2SNi460enNYVXbkv6jox8qHc7ld89ZqRucG5aUFeGIcf5iCMbBEmP+gbI3U8VLiuI
8atzDznl+JXmZABNqfM2tA0G89LEAjTqZK3zwp3ExbFISmoDjP8nA90o+ChpnQjW00wkTHU5uUHM
f+tLL8an5yWPFZNlTOt67ZMlajRqyCq3uEtvii426jiQRt7vpcXQD/8pdwELDozhVJpPDw+F+Yn3
0DQC6P+JSAeWYDgiUZ3rh2wEsuHq9Ph3rdCLpSoRYfSrdVce2NIPiXy8qY2hFb62g7OuQy4Jh1iN
pPDJIcegSBDZyYtYWqf8Ff22SV8By2WFoF0VjMCAkvCdpClRb8dmJ1OuwUi/0PMQAVVptFH1ZmRq
t3+Dlr9SZiXsMYxPfMgriU1DEj6Kc8pdE1bl/cGSzkU87uV8MMYoSj9mPiTAbapRh1e/zdYrAYvp
+2tuGdkEoOenA4Cgvss75UBaJYeWxle+uPcFr35Pp1O9mshpymKvxIoUjSQBC9UtVz5FThCBWvQg
jwdoE7bwhL2VNDbcpEL/hGnJwDYlGeyjjF69pLbyTk/B+20JIfLnxJgPuvQKNZ9cJMn8hjJxY+0y
nkrGHiGvlAw+SHD2khhdCn4r3KVFLKVLmwiataypPG9j7W+f4mHaVWr7IsPi3Gcreh1x3QTlRUrk
eqXeVJPJlXaic85kzVgXyZu6d5xMvKllscgyYj/u0gy8zeP46iRTx1WNWf/PmRIfWiC2nV3FGo0C
Gi53LkQS4/knYnXtz29pR72mC2h1Cnb2gHHXZdIoTHsSx25fD1zb14OyzOyIIR+DN9574maR7pUk
U5MgHX8vnFjMvl419SjLajPdxEW3xWJWAiBsOJYMDrR9G8Wb591Rq9hQAh+xLwWBEPOTK87b2ytS
lFDxce+XubeDCATXkuQZNDxU2yaZN2Fed4BNMab792i2o3j5YcAqy1v+DG8rEBQK6U1uVCVc8Pbh
PESE55PzqqdKCJyjme6Hy1Jh92bH9WejCm0Ev41wYM47GO308rE8DUOjgR0qvUtyGjCLHreY2325
wD204N1HqUUm3C2i0u4La/Hq6px+jHJd8JFk361tRpd4kBH0jIT8LYCoQy56wrYXOQL8WH+QIL03
I9Px5Hw/l1DIARuI2Wb4x31gHTYxM+n8XSq7oNKWIS5+aA91hWRv+60b40dWIZpuQdVovbdQayM1
6HL47s+eVeVn9PTGzelDulEOKb0a+Rhi5SiMbcl7drR0wqIxp7c94l9ONIgn0ahYcbTvaIdQKHiH
mbCNLKyNp4AG/5KIgCe3E1Ty5sHFKX7Q7Eg/N/xWi+ykxxr7g/B2nXNM2KL5pUUWk9Cs4OT8wYHt
+24rGtUTrMxF2BWQpJBEVUV6SV7cVgoiPlsy+XmLubX4EtXrW6wuXa5HI0zSyxRz3RRcVVgUBF5m
MZmDfNJwloc+C130XGNDbjyEMfFw+HfXEf7bzCDflSllBNh809fUYCswrO4v2ZaDfG+zMzG46DC4
mSbyY4rpf9y7AzqcIxFNa5bodIFfM5LXPZMXdasGwykm5+5CcNqyr3UfMe9oUPnuFce4pM5tapz+
t7bCa9zSssLn8/mIiFHWElogn5mATLU6o3nk+cg4oucDSPW/Bv19niP/hTv/nJ3szf4vl2QchFMc
DyBJwDs8hUx7I5q2YAsJIminzCkNgbPvHpUjt5ZsUS2l1hKLrpYsGewd2ggrl9DZB8/AHQnJN9Ty
l0GrLpH3HDPTqXcFyov2CYzow8VnK7GqyKHmGm+WZSGPaZeFhs9OOZw6PQvTlRYoMW+5riRvk5s6
6ACoHuEr32nVnRnKWDa5gju1jL6+evfBS9TUU3LGEdeKwfYbbaBYX9r7pxeDeRUx9whUpVDda8Yq
kECby4YO8qFRGPaL9xkmNtHcRhk1/a9zv6VyxhXV/oiuvyHrgbWk+NC8ARi/kIA1VGUfC5oT7UYW
M1fsmvZiZuvNKR6Uq2aDQ05nIZl+I+FDL+aKiCbRRiP4aP/KWzBIRqk6rm374nC23gIMdtzVm36d
7S8p5bSdg0S30cPw2U86vcingMXmqY8lH8tvifJlAmlFnYEhX6YHUABs3mq8JnNCceAhC2YVihk6
F13XghElpO7WB+T/H3/m7qoV1P1e5A6UrMBA1vjP6uiknGs6V4Oi96KiIuNu6EMM1YaeWH4Knoux
9z9bY1Yfdtv8vWRGnVqxpMWZLPD4R/lBIVRBS/TJjwJboOj/Foit147WmWe2OP3wshM9nthyW36q
M0MiPf+5cv8SrVXszTikrEHtiwHxffodIQRBX9+NsqJO71VM0nmxFUVKsNzYTVEvcTVtUEx0ElbJ
o2QZrk1LIb5BM9u+Jnsbt8PGWeSH3/n91OSfq2UxKFc1bxav+isczFOxn+qCThafwci9hcn4+/Jn
XlZtv1u/hLZkWFJ1vdw6WkOJkaYzHUXxCW6HfuTSt+NRAJfSlVSRUclZ7iQESAnYw47R1HjIocOO
JCGUmPvwEa5P3r8GfuANl0zpQ0LP+qsDx6/bsaZSOELBIiqeVL0yS53tXi8pm8wLU3GDXbR0UMqs
nQH3/oKuJsuP1N1qzNWKoHy5OOMaJfVq8DYU5mIenNMgOV6askALB7yP/vQ47QmR/DeC6RsJXMQ2
7uBcm9Bxq07yTCH0KpQ3i1PXZyG1CX733cKucsRgiZ5AQkyNDn+MST1blrpeBVcd3ovwXCLChG0X
zoJuF/ORqXtZbldAxe1ppFDGVTn031lE4j+QBh6z3W7Cj5MG64btHArMnwuTVOqhQfZnULXAUQwQ
pXtg/Poj2LszqdiEX58gjxGOAGtG2LWpzTEzx1nqPd//QyBTRLJVOza9HrWvnpaGWhHf1UEEt1+z
iMYkxJd1fKe1q7+LTOhyDVACtPNpq6ZZ4j6/7vTVnsW984qp/yo1utqUfWtf6PVbXlB5kmNYKctM
fDcBF4DfV47z3eqPngpC/4lPkEvNJ9ezCiTkX8pgTTU2mdnNmiy9JwliyINi2oR0V3BgEOxt+LmE
H6/5iE0lB7kIJujVmQnTyYHvvYbf/Jx8Jd8kUYN9jGonZdJ6dAIhpO6TmI7HkbQzlXtxiWM8LiO5
1Jfx9tKrEwYKNNsCVEh5JQgN4WNVWh39t0huE3HTYTYUN5LZPcYHaXWJ2jLlKolshGWfBiIeoIcp
V3qiPT7rGTA08wFv0uCQDb537b1jhX8+rTtMqqd1RpZJ7Gxc0vrcdeCBcsPaK9M4H5SaSJ1FDnmh
kw5F+QpPRCkTWXp6bcsI+KhsJk1+1tdnLTwATwlObEyb7xSGzp8B+XA9hPssChDj5yCmJcnwlOFJ
1VQKPjB/XBn7Wu/NycGQBhn897bwFeasGwWT9E+144nCqa7TDa0xOmaH9g/5RGYi4IGUwi+OMdz3
xWbLKJxBSEhiUF3NjGbl44j1wJXPD2E/8V0pqAnN1TsWYtkrXLQguutGn4X9W1Mfa9p95N3z/qVj
MSeQw1tjJgRM00hRkTkb81Q551eNT79fvnZ7Vz5sNbr25a4k2QFPDvHi7VVvvrFQK/QDGyLBDZQo
Q9keKS52WTyHBmZz3BrcTApkKvfeelGVfIps5736BNwBJ5WWyQi9D/LePIJf3oxzCcHjwE7Uk4eS
UF6qXOe8qeqaWlzn+mMNCurPuIKWalB/rUrc6HKoSkNrzoDWAMYNdwnFhLySUIgTuhlI4TTyg91P
QmzLfx3sbXxxDkmoDNq0s/DodaQ17/4r/sxoL4d0
`protect end_protected
