-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
B8wshhATc0sz+Mkg23KsiBMq3WHatBELFfEMEMXBDpod2Ng2J6tLjVjA/lsjc5yd66zGKeyw+ntn
ztCp+ESHTbclFN8mKgRzp75NocK3PRrxpKsAMDryRUIqUhiFOv1e/2hijkvSSnei2e/VIdVuSmiD
3Fv5Tj53U7ZgN+2wpftsOqYq1Ffkqw7hkXmHAsGJcKJjBIcGe6hmcx/AT7c+GvieMkpOkihOr/Q9
n/Z2Dq0q0j0uHZS+xxeG6f7c+x/lJDQKifEqajg+bVsgqAe3dVgi3jqVVfPZtysyxZTmyGofESxw
2gC1fwXkQ+9w70R3s0gNkHSNTE5so8/BZtB+Ug==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10336)
`protect data_block
68oAhuNaQXyJ8+DoxIPehcRax4VMiMzXi9FIBh2fByo3QKvM/cohMJIQUau/GC0Cq5kh/L4IGta5
v4v5IR9KfJjxSpvf0ti2gN+/Lv0MaU94bwWbyJfjS6N4M2PdzLdbXf0PoVwHTaHPolRvJkvSZ4eS
GpPEG3fXxTxHebW8LLBCCCFp7vDHiNUqXE19TeCdqWv7n6q9++fOpGwCEnHf1SP7GR68V46Dvndp
ktYEoC38U/7NrND4FBryIjfsww+Ykk1hV6szDMOfPwrH2n6YApNa+d+MwohapaAt66pf0jS/H4Mm
aMTxyCyZMPoeisxXldnQ9uz3sKVJ4TzH/OXjZCNudnMDgp9ECjslXMXh9/C/a4wphyDvpl8gvejX
W2pXn6NgSIwXIMUuzemKcFTOLVtdzVfMxLNXf9gwgsd/EL1qxZ5GCEavtQEGkUBRh/GaJE8y71DM
cpwuYZPgHaXRnHINwwuwIplTyMsqnnUh9Z7ckSX8eua5J43yeEEtvBMxI76kcincW1RbukOgkcdS
Ts8lrEd9Gt7vlC7wyH5Ed+QXb4KNd2g8K92jPDN5PwdS+sWcMfW6odO7hRctWFgdPkaEvhpB3CLg
z5E6XoBh+ZVjen/AbyirIu9fuRPZAaH0Qb9rBuv3Wvbov+1az2GqI5KxibKne4M6rLaFfnnvRYQW
h1o92KW+s2JzWz4Yg2QyvN6pgokPhlXNq/ADr6tbe6Lc6mbmsGsEHC2iXgXeIm+7VD/T01lQprLp
ZkZL1W5GaFAyakCqk5p3wBjIl9nk8sKLgo3DFL4jymjDqGFwHawduNFqVFasko65KSMUZRvpWma6
DrUfny8IodHaKcC9paWIw53pNY5F4GPV2yRKPKARxVvYqxlfOw5NSdh998ihbsoTO0n9KWDcimxY
IfxzF40H16entyDKBXyTKwVrHbIIA1xlEOlRmGMDxmYgYDxILgviv8jy1ax9CMjY/EwSd6A+egLq
R92y/7rV5qX9/O1AIdJFJu/WBe8C8WrUdLEYKKQfs7yMkJlQA9/HshrRaAhn03WnBnk/y49EOmJ+
N4fGiIugk0A0yRX49KPN2cRUgGaJZux3bF26v9w5HToA+rZfYq1Zv+ifSN8b3zKQKLM5VzEz/Bo7
682BpuHOvMF+7FLoImfWn2sOjzim+viH0wRtwoeyU2qwVp1Y4xutymzECWx90ZXtjM7RTbo48Rhz
73Ztlma2aCssGcgnic3MooF/X7ycAjndWMtOFR9bHRIlxbkFHOCPdudK/0kGlLf4UL9oJvUC9/iw
xn1Ka1ovOWdg1PyrESQDP1uI5QJJJQoovke260V7Eaeh3YXK7rNET4dS3Mn1Ca/glFxbJBxrXdg4
r9Lm/il/1PNX1E2SR+juxgSo25ZYovmSYdlWcoxMEDTVn5JcA/WTWgMoXC72eKvdGl1G6ILwTnrt
tLiYYv2kejSBjcoD51+A4cdmQvUeR/gELuF5jAbD9wn+vEb6Fq1v4Qq5ilcfILZOZdVHDuzbszKU
2yudZHOKPH+dIq+jxb7fOzM9k03HstIxSTymkw0JtIIHGBvK6gr+35lfSfOB0URepBQkzFMlWWSm
BkkLVzkWZFT+n+FACG8vb6rpwhCColvgH7GYvRvUcmiMTRPVFVPC/htB++n/fCk4depIA3cuothT
7roWulB3TBbM+A0FYUWGKkXG0ooPu3tTVukAELWTapJYpHYybV/At6QDNSuF387E3FtxSa8qHefx
tdnyOX+qsOwPb5Ms8lYJhsSA7zmUnSxJqahFxO0uYlxDypVh5eE3OoH75uAUNgePkdpV8dZnZ/bA
UK+C12O6UKmik79EU5mcpqK9cLlQ352uDfhaM7n3AZi3GCmVOnZjedAHvJ6EmnVFG4gvbPlayWMH
4tSge9+vL5v536C8uZxUmkhfCRMvqYCQbzc5P9+vftDNOFNsDfV3HiHK82a41xND6Q+4+djoNgDo
FwciTodtvYJaJZsqihUqlzRrbOsNbeOBIaY/LySTVEFSfVagBfrFyio2jo8ryrLPU3qbXqPe+7k2
2kkGwqcRot63TB8lRCRmyXhsnNYt5niiQ9ikYJ+uxn93PVUUdEhpWTNqsKykn1YOeqXB8WH3h4su
wAYe2OlHkzv0VNqoHcPeDLkTA8aT1NjBHnfQ5Xt0vvTlzvWhA09ssBklyXKMDWSibLuYQTG/yERP
pzMkK+cJLfeucLR3sGtna2M1pvX00kUmC2+FmnXNK85QU7MYojHxUJm4QXf/WG+71YZTnEjAjfYT
AK8lYNL5jj0jiZS+iu3t5nk+a3hjAIyz7g9kLyBNuauwevka6HW7uidwM1iK/CJ9M6pEwys9v9HG
srWlSndE8SJGK8jxnTo1P7REQ9F+OVbweETPP9aKjfeK3lkwqzXJzXJle61UhzrUAAdOC3KUXfyY
d8HIRGZKBpVv1TTvUHrzDsL0G8YJRAYRI1Jfw72GkuvueEmYhYFGyRmFdls//vOreYYrr4WWhtAH
X7UAbFqR+Z6+DY61SIeFGbteqQkdBkv6XHx7otSAYk3CaLG+ycQZSyYsJZjseIxyBeFyVV4a1zpO
wauJ7iFERceWvEB0pAXpUIINkgSAFhLR+0gQSa5VxZfxadUr3aisEVKFjgc+ueDqB5Ef+EmHMCeF
VUH1ZRy0ffvYY13YbJxtL4M2DEC6weT5J2lJZbRicbeTFrn9LM+q1TBDusvzva7+UPhRphWEkEQt
lwMUL3yiW2xR0Vbeh72S+T7MwnkZTkV8rreUZZEg3QmqxapLDn1JDoiyyCS8rE4BxalXwsRgk7mB
o+TAE41f3ExvHS5PBYuQaLo71QhtIOIDF3wp+jU5lsyMxzwTXkWVhwpXtXriWuQvyIg88lbytWBe
FsC5sidZLCraGW+8Zge0cc//y+N+OngKvhY+8ptqnNuVlqhtksMuoyrAItAFSh/7KqNcU0s6vvbw
Eg+boQDIPnRaqE5nyxS6ipC+XQXJHIZG1z2S7LyRDlQd+zLS1xNTQJqrkn/28gr/+qnlxPYkMGQM
qXQWSbHcmbfmjBqAS5tc3a51K2W+UuI3U/cm+YgwWyD7gJ3GkPPW+bKWJerfbdT+HuP3BqBwVxNZ
oKgTpzUbTj4M1XhWecGJI6kAja/7I2NI1K6Dio8BhgkbR0q0lwPDhWvmSUM2TTz7ss+MUly3Nljt
IwoGqOCSwMRZi7F4bF2BGjaPrnSZ71DMlRy1MCJ5SYAhcyB1QI9NE5mjH2AEzljd1bLraGET8Gj0
l3hhMLWAVx6GlC88/bzM4Y7OMnpgvPNaQ9Zu+GekgPD+FmxZDA/x4DnxTfEgRDkpf5gaMtTUnOmY
dzKY0iF0YMt3ZgrDyRJbSzrA4P3Yqm2kFFSBLaLkhjTvWqWll552nlUSDjp9YmiQZrhWeGmBvXjI
aa6+DJ/Usdw1X29ayJfXsm5j8pOqsM3RES8JXplW79SXL7Q80Fkkx0RgWaS8fZ9cxjCcQ2cKsZqZ
FQmeVwhSYXwSjFQ2yoFfdbgS3CbW00EgXBpewA0cwKG4+dO4rZGT+/mNCQKARSRYuGg7xRFNLMJu
uE1L93rPWoevIyZPNYAuJXOmcvTIKyvDkYmgBg05/HAGQgj6lhz5lzeYJynkwMmSnwEcVld7u1PP
EBkum1H1YzSxsBs4iK8hFvHpaIxqa4bbbqLbpb7uQJjCls1p1+MuUlK36UMbGT/88s9rN58Ft0q8
87hVux9tEgxSgZAMGWbMJsN4QdU9ncvpEvFTU3JgOmAR0WGXWgu1eSt9eWfylZIn81vK1t7Xn8Tu
iT+P49XVYRAvpsCQ7DOAWs1LklZNimiLyLH5hlZIzluJvANXf5H5j75/pulAcYBiXOMLRBny7w+k
vgdNTKamiquemGEQGnJE+0UfgG/T3MTEZOaf/Z5l0Bjv60pu2cf+kTI0AKDxlfyUuvDxKQj73EJh
cmdzYodBzReIhyDQFX+4jsv/SyIFCgGriwQNnZpIkv1IsfXJVyKBZkOZTMb5sUQi+JLAJy3As/ry
mpIUu6KAHOlLVDm7DhAR0mxn8BNPE4ZeZui+QWNszjSlt5LCwNNUvsVdcO3VzsOr7/BH/exFjxlA
PaiDOCO0RoXMmH3SHfp7iIBah3aqHfwEm8plnt9VCA8g1SwB7piL3innnNhzBZtqDCjeaOkhNTJP
8maUex6vQ2yCpdwUmNWFlmh47SlRlBcK/A9HQ4Dj2V1TM64ubTFS/4NKcOmfWRQvnTpNSJpXbD1g
qeKDt1q5Hzw7L/TkMvxLewfDrNZ7f6pvD+a58HWOwg/ih3hDZxph8UsaF7vfSesnANiD+ptwPFRG
a/QnutXoFHj61h9uLsUVN6k0FcUFu9QvPXAp+2uXiLL4t1IVJeNlvGvCLC19mFBVnYM097nU04/M
18PFrvH+zzoiigAZLC8kGSNq/wPzb4ZLkPCW0d/W7hIRhr0tGXWo+eUYkZCs3dpLz2bWC1D9AdZZ
NT2+wJQD8v6wL5T53GfTUG/Uy3W1TMKv4w1qhhv6bkuw3e2UfjWMMiLpNRbnfVCq/mRIC8w7HgFx
VeRF9mod2mh6DL8EyXcEuBZjlJZ/z4UBuOPn98MfM150UucJfsoZlF982ollOUVkCCgRoEF6jhT1
wOuy0XFPZhPnybt0mvNqGa4YTGqJq3NfoQxNGTqbjE7DAK85pfjO2jyBqgMBb1d3KRgEGFfSyltW
GMXWXEQVO9YBp71qf90CQOIGePrnDY+F90mIqg5/53taskg5M2ZotCYorEY4ZHUjs96VZSRUiUPI
x99ht4EFxBBUjWdkL7mUPzowUtf1aTzMCPfOOHZf1t/7ufM4LK9EXzO7anfCzuWCu6dlKKBg4M9U
QQzzXPTzSw4zlzXOMRS2V4hyJOoxDcpKw6UOfPIkH+7JHSGpOmg0VmIB2RwjgiUqrUPE0xmNY7jT
hRXAsRty5EBL7P1t1nWJNXVESeV74qNsmsjXGKUw+sQ7vXE6omh2y4NXXjAsbGKzCUX2bve685tQ
fHT8nk1rh3EPTA3gVBgxEZzzGktTTYaUa7IjCTyEMaxzL26RJwcFP2MebiclWgBN5WK/zSW4c8H+
0OPQ6blULmqYUASUuJ+nn8uAFCso06rZ966irfqHzk7oPwhkEBrjp3yzE6VB9vsaB0cr53CZ3zJl
8wdiu/Th9awUiq177GXGYVADktBJFQNvqXGAAs8a+Oep0xu++jn9E1S1ETDhCY2ViQz0HG0nvvb+
CshinkbuC8aJ91lACRGkgpm57ENvxZA0pqh1OnvP67IruVK17bUwXVg+CHcDldwFzPIqUTWtzjo5
9D76yGe1MtDy5tJTDGD4HdbS7qVH+/APFLks+gB8WCTo4GrmxZj6HGkca9R3bipsZeCQhU/N8r3l
re6pOHVFHBti8eFGARhjLZa8qyBpD5SzO3c2ebYhvSW37TXwk7nBb/uoZJJeNkPmoGEIzt2tdFqb
2+V27W2/oJI+OUZ/1m3AsyIj15fdw/bb1gjWtxpuCyg5yuQeNWjNeUiPVf/y2c8vWBXaV1mJlQ6v
wIVMfSaajdXhtmy1Nbsgt2TCkDnmtGyMytHlmKHipYW26xgCQ224BXcrCLgfsq6f3U+Xo5p0y9My
cIyDsUkX6+6FqqXrieen3o5cJRC2TiWkXTzorybkPuw8BPnDPFpVJ6fho2B3xfJVHHiKKICi8/Sr
afQTf09ePmUnaSM0Ej+PJnPa/ySk4qtUIl4K5YFTGSKInhzvV0wdp9OWZiX4Px9dlUENHM3XwXWm
6b5LFoLAeyEUMf+h0gvpdKaC/d9ktyB4klHhtfS/mMFNxmmetumeI72DIr7KvECSZ+/t9iXkrm6k
Wu+0kuZwQ8UwGfcTD7ryk90Gv6G4rj7rO90JfPZvCiwOMWvjfFb4kyiDTKR0Urf++eI+iQhJeW5Q
mpKJzHy307qeU3HpciCzT/ZthEQ8v9XqjJm0hWJD7xpcQi1F0gu0R3Pb2RikCj5LiDD/fhkWCoLL
VloL4NYyM291r4mFjpQK/Bc9OzoYcvbMhzgplgCeqG581nRSx138EK31bi+EEFr8CQTn6EmpbWsU
3wOKiH+iOAIv5EGT9mdIZCBVBnwoO4Lk5mzG2l5JvZ8uJ5zAJozJgRrrVDWmuMZEtH+phdH672BJ
6Z32qKgYRn/sVvI3YfTr+LGnqs0ibNTMQY5twbnASDX25TBrlkCJA/nNbam79fEiV8YRQ1eQxFhw
uB+ODmHSpvxduUKuM+ESdo5hmAKzEXfwojPu5uoOxq7Kh0kvx2Qv2ihTKVR0TeODHlFNsPM4Gk/a
LP7bL8ElbaWJvzSkCEKRRN4HsSWuISby99q+hSBUkznJcIMWMmXnRaIU6RbcgyjFwJoBFB+eklTq
0xjuLkcCXjHuWkOSoBGOim/SraHQodMBRBqtbMP1AIq+HcEaq5CBy3Q7awa5TnXv48mdZxXgnkUT
5A8K2jJrbF5VBTV2/dfIa+CH6UTtLFHyoltbgTnOWw1yxM8E7oyrrWKwoiPo+QX7S3835XLzOL3O
i5ZkOaSwgK25OArUX/O3uhHvUtwpQJWnCJjTtP6vEhkWLRIAradL55MgxwigmdTY2yZphR7yR1Vr
UglVuji00MiXwn2HpX7lSol6rsVYC6NC52v+pOtzAOA5VbKCk0l6+58gNQ+loHPoCFSRR8gHCLjD
HkS09ExbtCGvQKbbVgQZ9KVsUT1dnWYE7uEVmyl/cXfpgb3T6rcfpI+bpMeE9Pj0iY+A3Tdezl7e
Ob1uOEzBddVQaw1agbPAO3IwspV8MThScZe16NYaabgDgaX0d4Jq4Y7fY5NLl2bWyY3+4UBFpe6/
0ZheQPoQeqkfj9fse5sd8qjcMgjR5yurIYLBaSVCbyWlNn5EK/l2yPUOueBw9z6166WKZcRND7+F
gxQRMOnIJSszAuOl7C2Ew8sZzdGWbQcrJpTiVNjUz/SdObNqbiPS+yLX/wijgC2aHDHo2Vd0SOVq
3UYm1cdY6ws0ZZV4zT0Rl+Z0oIV+q/awWt1rj+FXZAksSDXPGcBK4j8SMGBg6qmg+a3oSh5o6lps
ZYw0enuD4lvZ5ldmF65EeLAimCJXFDmdOP8DIC51/MieL7hUbIukTHgZxmekLk+IdmBLBl/E3uNA
ANJwVPPTtBFbtm6tPn8E91nYQqUcCM+V1ykQMdqIGI3N0Z7IY4LCNRhlrewlYRY0J6YW4RllK59G
OSNzTgQOy+WaV6LDM6p2fx2j5U6hMwffx8cC9eXpTqt5RXdFPQ190uK3Y58DGxabocTCOx77a0Ex
dPG3ZmyQMla8HIwwU1ExUpcdONIfemU3BYQg3j6c2gRx81A6J7donytedwm6gZQIfkuPI3dMIQ0e
52fm6KcfnCn04S2sev0RWmSflKEYvWB9ccaYNBFdeEcy7317uLnw794HinFQD38sM2UU1Yq/us9k
1EJBxAopu7MEG2TpcTYlz9z8cgB0ZKWK6HbW97UXcHQyPq4pIjbgPdz5GrPZf4l2ugCBVBGjPhzf
ymIXuRw7RtkzlxjHvX2samhNR6QTBU86ab1xFfzuB4KLv7yssDPv0gLe3XRUU1tR8+NSqWEIMRKs
1JjB0YAqcYMK1K1nry0X1lXSg00tymqlu10wgqj8KQtpLaEJHKP2RUvp0i71udn+N1D0KUGk3Pv2
ZbAKehoFeoUwThDgvZEOe2TUMCsUuPAAJx1u894IKtAPJVS6eBAp72dVkyu/lV7efNNduFPTEcGy
HeHKk9Oau2TEHBLIEjW7HrhwTd3jDeFoAhq8UAO3L6oNGJ6LkO5/I6aZE67Na9G+jCmp/iTN9sKI
V+CcYY4TSotpmxNevD49EucpdkuN6kbj+P1MhIe8mAlXmtB+1SxTs9Yy3zl4FAq0582gh3aL1eBL
7bLHcOSyVxt8VuaeuQA0KMB+60euP8SpSx08HyyPGVqSOs9oRTkldtKmbsl+BiWwa37ocyZTTHoZ
5KzhxlxNBsWgLctNk8HiZy/FelzUQ3S6DL7VH/5vRR+VAw/HV2QVuE/mC6JxsRTTe3TRT++6nnm+
KFYef2LyLIpNRrfQOh/tWUJIz/zaJxv6XahMa9577OHEDk9ty6217UuB/uXH9yPHheQVelxLh+Cz
4ZEBI/afl5/aw57n2f4CTSoJJSEvHIFpM3wEf0bEc789c2CQ7/ObZJrIaf+7yoONJB9J3I24kokw
wxB3Dyhyk6kNvibAlInR1XfpGGVbJKybMiYXA47XUv/362217S74wtKbGOd8wSkb8242urMWYSXM
e36UwuIrPdOVPfToAbjcrGGVAon/C0MNHk8XaoBG+ZqK0W0VE9UgMR2/g/HiIR4Nh4sqGG+C5zWu
SvmqOad6lJahhQn3cEJPqdJY91CDJhdAfSI0eU8uGGiXYP3T6JRuPKI8pHFomhHPF6vei7Cg9dr9
Vl9lDZbx80UhvqKL13/uB/InT0/is9Yd72zxmdPGhLFnNwc1ck061r0V2HMDlQWAEBDxLrmEowbn
w78sReYgE/Vsepk9o4VH7iv1OKHOBCc24i8p7Jce9HUXheMohKDBcn5dbfzyixO5rVivTFqkGhKf
C35LMdK137y5XgnsvV2+aQpQPRr2ojiHWOoqShGSFddxchk+eK5Bbo3ezDPatWKLpO6oZoBh026P
lliLAl2wwtRY6vLUpiNVUArRdZd110do0d4DpfjARfFi7ja/t4Lm84laKuLl36t0uCZVIh568E3K
IQ6TQHAFYFsHY0YuYozKy6NLoym0B4AUTJ1KSkbKxEv0T9d0dOomwXJfFMOxqDYK8aVkjx+OdRbG
f1AV1Xp+6UfcRwWHqcBkxDiCTH20dDsoz72ALL/Cvwy0F3mpHNZFmTh8K3gR0k6q5FBFwV3/iBSF
tZMHS0Dt9eQPlw+eMUY8AfjXjuFpHSS81EPUePlxTueWLuFt9xyd5Rt3E74Jvd3cvL+zEuzohy/R
5b+CNZbJCejikv4+wnOFEKQvC/ATzEPT1KXs3hBDaX9pNPl/q+EGfKfqpDYcivqb0ivEbeAoHq3o
HucERmk9tk/jr/uUEMk3gZOIvptwODgDZyLMUNJOxCjRTIndC2uDp1Wcz8VC3cn1QVXfsiKin3oy
MlBRF26PYK4hLg5HOz5rerk/b9fl2yTOWAZpeJIQcFN/ZmzEprxgMI46TW+WmnoWYld3i5gV/mL/
gJ4SRGbgeqMM5mVTPuMpeoi/2rNTi7Shvq8PGt4fh1YrE7TS8G1PUvFGkydJI4K/VCOSK7eoKEd2
G2qyQjp0V7XqGERAMH0YpgQ5vRXQrUn0dWcM9kc+uUc0FtdhVFYzLUASZ8B6+VwAemJtyNIevao6
WZesM9j/o+zHN4tg5F1jFP0y2cUUFLb6V1OjwVtiZMAmb/cTQ9660bJ5QS6qiodtJ8B4RnMv5BOs
FURxGzYrfbwWLJNvE9JLa/+qIMKeRG6oj632QX/k5rZfTaYS4CNcNH5ghv2EafjK8c6U2qOLgPVD
kR55frsUvlp1QUkj09XP4ES/ooJTNSn3kTfSp4uItNK935hG5s2mhZWf05jSIak0MqJ2xruqMTp7
9reubOpujWg8TgSdQ/VrM8KNzq/4UlPX3WApkRF6NVSP/ASPI3eLn04oVOv24qkJ9oA5Jhd0uGza
5htLS9PFK55SMdJUo54i8fI+sWHS3WrWVZ0jGjEK1akKV4huc+pld2x+a3BqqUjQaGyOzzwQxkQe
LnV4VbOkZkf3MImcqZi7F397h7fcBV8nJcuL7JZg+Xfu4Mbn6Bcw6Mjlo6pHpIUsLQIY0oAR6xHV
C/MNtdtH2OW5UTkMheT66IU27MkBIATjBs8CvBfL6okdu5/+Tb3/wzEE8N1DeWaCj0+77zbW/ivA
Z0MbD7424TFztKexiw3Ei5Fk/PsNCVo5cv2gqixkuMKEh6IxVXOEuLIsFPQyyQowlJ3jZxnFBVSR
PeNKUWnUz3NsKkKvqVgSC1FmqSiOM8DvJKzSk7nAa5yX1ge89NboHpKiEfPf2Y15zdE7PPJbHLDj
3PNjUXQwg/Y0JlZDc2bdzxC4F3qZrIYBE0Xdhhd8d3IwLQAF/ICQ8iXZQ/cHZEe1nFtLIALvEG0C
x1l4keCm1p2pnLFKxRiHgswtn0JfSeR0cDSKyh0BM1y5MYMB14el5aRObQi2nIbzd5Ccn/YQE5d8
QgHicr5IiCyJoeZA8VgGAuhv3031ewqlvZYKj4/fifdspoe9YBrDojqgy6kqm3OENI4r2dK9fdki
B0xq3abv3bXMD1WMgRe1qUjvgt8Z1sv0GGCwS6GtWdH3xxvVY6J7fSYh8/VXaVoPg2vq+pUz5D7B
Bvg7cb+sHmAqrp99ftuYZjVyFQ9sruxiRzLWqHPSbUm9nITAQgoSReAK/SPQww14P+AVH5O0QdaV
bSJkeIFX5FQdXn5aNU0gYFyw3YYVXtU/bwXVXPdSYgKo4qNYXsa0gb4yAP9xY3o0lLYHYYO5Mpzc
0dkQ3qXrk5SZIs6lWRMNWQfHNsFuM5yNn1VMRtvdRQXrHEfNGBAbxP5b5dgTJOp0gsTNviwKmOLZ
gfHRFilGCNKSxBAdif/pl4U5ahyXd4a7XrDYNja0RykYxuu0CHNpkvPZvYyfZBwMSM/3+nroGRHG
/Euax91fzMfrkGLZGfRUOnxoFUWVT3710TWPHtoQF0NkW9pz3S4n4MTBU89dLqhXkjWOnchqTLf9
RqlCbWXorpymq50p/JYSKKgsfM9cJA4Ftjmd4UySrtWw94HXSriSQrK/5PH1znL3vSlQd4PSm7Rd
IKwD7dRYH9azHw+t3NQ3RgvJ9bjHTZZuZpf6NBvJ304HZ9T80XMlzqPk/4mHkm2zqifrtxvEQEp2
2++aHlqNw0jXojavIpyA+fnSvoofHichwyBFOcVtTuqLtIzbp7lLoOR8ymcQ7+vMzBqfAJR0y14U
PVzmVwAwd8bRvn3he61OSIsOJ93eYiy8fmsZ6GOrWWq1d+OQXlcqm00yQ+3lza0rJ4BJr0/RBR7A
wNbqvT66BCrwAlCPk5/9p4MkWTcuuGk1/34f8WgcxjdyrPGinWDcypDqU+NUuMUMFHa8YrwkLvtJ
v02F3wB9d+PLUPcxTt6YIlfRmDt33/OA0AfI+0PX6l2tQ/iJBebG0kr7ZE+uNuWIJ2TcjHYAe4li
DRK9hutV3g4tErAbLb+Xl6BzgEQvTqA4o8eGjOk7l4QR+0x6TlAXrcnjYa5OoT7OqJkuS0SWhJ1h
6MxRLHyAXPlx4PPlg02/T5Wl+9dbCsjIXRoE84v16ByG7My/Y+7E/BQZccp+OhGr+WOEC5Sj63dI
pMNzkL4KeGvzTVftRVoL2eHaY46dHawlegGepD6g3wAIAgdxIFT5Ne6lobSrz1UWdWy6fVSDqMsE
NrABza2VQJhXx8TtVnqyQAMz+TXnp4qpwq2JdPcpfD6iKUNA7PhHc51q9SQ3AwjAGmLEVJibLgv3
Y8QR/PxhzFoAOLa19xTiZnbYx8kb8PEapwFSfCNa/vs+N2tiYFUYf7mNqu1xEkRrkFOJHDs2GGtK
kGSNDLETW/LARfSSvrPILC+/TWNhY74rcGmn5YL/SLtGIKqXkscWfJO+VRq0V6QR+Jw5g0vtDkSO
Pd+hveD8q2b0DHzqJrLcHOxdG0QncAHT8rzfrvIEVaPsEXUPZI1tQ143/wCvJVaBt0jyH0N5KHWv
cKzk+7KfSVh9LKxicQYSI84QKfHTUhpDe9ITB1WLkSzfforTiS7b4u0nzDKeUW286e5ExbKCpueU
2IH5GF9BfMDYDvG5YZKtff66FYYhZHJi8tZUmg9FuBlDDzQ2iQVqc5Yk4yVMv4zsZ80Vmgn217FN
vmPr1HE+Kva/gLgA+BgjIHVo9OnH7mNfSR6dl47bWN/jGptlacosqXqZig7t8ST1HDjvawRkI4ne
4YuquxRCqIJMn64yi0rB5PKzBBhWYUiQ021ak6HcfZ8jFKRTHKKs5Mko+xiRk00DMTXzOg92hTEI
eUgPCNx69gX8HVabMeLtOh+I5TO36UeXYrApyLKwZAKdmaAgBErjCnlSQWBawhTyfdSOLsCJ/FAu
C2s02IAYR3ZJUHhlU8xj/S9bA0fEUs1hDtWrBfL4MtO+PfFhPd+XByQp24WRmFX0TE9eAnb4hawu
SGW5oneGILFSY7LNgKIjSCjI6o2hxa4OZMciFhqhzYcuqOW6NKkBNuJyOFLruuFGFnrcjDryq0fG
WhtLNjXQ9+6BPilP/PYBcdRXnQ9BsdIAN1c1A+7x7TmzHfMW6JynrSiCru7v3eKtLOtfBeEaWQ8i
b2mRFiWy4dyaBvBmtUt58O+RMyOPasuxzrxneIs2qts58dWrZShfk1MRmsE+Q1C8WOy5aFT51OZ4
YNRzrCjTAauOSa22on3Tijfqs6AbTWxb0yau4BgvmjVs1yJstTyFjM+cXTs88b8+JHXhQHjc1GG1
hVQPUfGa2ITi7RgdzfELUMN4oGB6btfNFKLJUzw8BVJkKON+x/V1lUa1uhbXEqmzC7PXIPu/MAUx
zG2zpKcUloJLec69CGx596EdfXDIByrHDgpg2rMl4sn7+r72/xrKJhxD0SR9EjmJr0zlkgkQYguv
26H7zvLxllBg3ZnzwqBz8FCruu6mRcvFzlXIMk/zDY2u5YU2CU0octDmHCx0uHTFx4r6WeV3wy2y
QoJgberfXsjEwXJSNqXIUeFuRjvjEerk+Y0z98Z8uSQFqNueIos+6v3qoPREHr0zh/Nks8C0frtD
kr/wLXSktlSLg0dWPKJtIuPk72zJeBpjz5DPFC2p7dmhNPw6IpJ57c5f1BudbuzbyUsdcsrMOASo
1N3mCpPEo6SUYcbrAO+arkdIeRSqioFpkdODVo2uhIBq5wXdoduR53rOhjIDscbfYFcEopYIPRy5
wedmEBCgCA5mZQ7ZT4lHrXB+IHPHujf6+I7iZwC+exNWZDrlft+epkcK0T3wCJXi5utFlBYL5RXV
nrQouf6Jp9pIGRKhBlz88On4Hslocff4l+ZzoM6uhgtOHdbhkdVZxkoKEwAgxszqIGcs8xuhEkHf
eUe2K9a4BY1FmaNdqCZTUhVMmzMc9lycRTcfZytrsfKFdsQFlq1IQMmb1m0VARQtwTvlysUtY/va
ip3SPYVicm7y3MjaSRH11YyWwlsfNn06qnaRnlCVLcvT7aF2PlTbRJPI/8ijqQeQLSP8kdspQGUw
Rp8N1XlLMyuVAFISIgjKTmZv2AOq5feJ9aY8JGyIssCalQxo3wJuO23ya5UTBCAq/rQDH2W5ffvd
CN2nXn1VTDT8Trh4We2MIshtkvtF+PuD3ytfW4uHuLzvEbQIoQXyJgvRkRCGxNdgYjYflI2B7A87
PSaeld/R5e3A8INyZkjepxDhvmoxnpITNaz8oEYx2gS40Xot+4YDdDngt5/P9aS+o3ZRpAqWMLct
/FuHqzPAx+LYjgZqWRdthgqbodXVsuEKCyp4g8bQGclmS+fjJfGCA8D3yVHlZ9mSrmTLRrwwlu91
NZG6kfbhaZ3gW/mpUgtq7weh/CNLxqsRsVoAK036WIdgb0+sAk8no/sWgdoMljqWvmeTjK9WDnPZ
q/XWNimP1uw3uru+FiZJPfoCU4RLlR/py+J6WawtAsRNuJstzXvyI6RBiaRASpAVYFoSaJ+pOA93
V9y7k9hY6MnWP3DF8HArZ9YtVeKlo2av9lTkePOWs98WGzYTbfjlsqIFE+xniNXlEOMEm7Sk2G20
cue+bmT3w86u3aGM3TgUZbSu6w==
`protect end_protected
