-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
y+PjuaQvmgd8e3X1676Mtwv3bFYwnYsaw8b0Z7QzjDkhR7mlkC3CXYfwv9bic0PYIR4kyfVdId5t
aL+hNpONT/exCjELX3+zYVQiCT7QRrFqhYhtZh1bWd5vdN8eC2VninzhGPYl0A2oq5itsheHhJpA
r2fS5huVDXlorHzP/JZKCBkI+hSoJ1r/qTbhRqf5qBsUdRCpzLtvaeu6YkcqdGUkF4d2neY0NFIG
R8UzKhLWbUrI6rGwkeULCNV1aNeovPhgiBDBZ1/Aw1xgQ77CWIahDqVMAorBoXk1X90r35LBcd9+
v1lBiW+wyOMrOVHII8MkhiYp1uwSg0ucnH7khw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9712)
`protect data_block
KWoxMMyVsz8+CohdFGr1g90VUO+5ghysb8PocbkHi6r0mBhVJEKzG4iU8KQCiTZ0FdSQGOyUcYrg
OknX8SjMX4om6GOFKaU0eDhUBXKijA9uv6grttdOvN+fJ2DtjrneOntMUnAQjxgkQp+PZl0Cd6O4
vF+zXQHBv5IQ7DDdOGd513IT/y1A17o0lZ6y3hFTHPobzgCwknWqJCKyIpTmuvNJ5VTNyYjmSQQe
OW7yH4cjfwF6id8qP5MVGO7m2lrXgU9t7hMXfdTPvnrCpV9DCrDrEFddWKJHJrov0uhsI2nTEgBk
RM9fl3yFJeyxrHFFNtEtQc5YZ4TZ7c2Atid4SBbf23XA5d1liYHGKXIHI/XdP94F9YHex0Zrdk9x
ya956gkyXn0KDclKOLwGQeBkqIKiaW9R64pII32GbykM/6mW9SGV5ryKtxVJ4SEh8+JBv9HlsMgN
hkH8XwjBw4qOcVA7oJIbCSkN1RKMeLKffa1RAPighHWfOisfGSJvYkRyHe5m84rUqdpWkW9hjXg+
ZWH22nvBYtAH3lyCPOTH0/0Yq8riAfvx8FOtKS2jFCKZ95BGV8gAa+PM/xr5uVaUfY8hkmi6PzbH
05wfErvnsOHxrraedHGaOSK8VcMU6DfnFKkstUU+7uWTd4EXDmPIYAnJkKx7D9YK+g/PLRs48gVc
d34wqiDx8dxYULIb4jPUGxukrhWI0qHhgAj39YlYwEHVLCylvjbZqfmUqGtsLv04rV12/VJV92YX
u/+FPIKFOpJxGFxlWEe90wSXQmnJBNktYdQZ1v2wTPRWcHERyAIc5nH9zzUDTmAuBaJHmeDgBPEv
2bDO9FzcjeLfDlY15D8EzmZj7guxqJAXTsyccRnYSWbkehYCg5j2GPSm9X9zC250HNfnEAscy0Gd
R1VMuS4YaV7v2Jl7u8WA6lcNEVXCGCLWxtPie76YVBxNdHzTm1sirguokoBARZaXsHMkmH25fkNf
lN4/OH7hgcngHxa1kROYGZd7UVCoMry1ymEwHu5VV56LtJduoMjOGFkFpjaprBM9polJ0LgHxKo1
4n7AteODWTmfNNllYT4GQToiLnaBunYPE7aL2lD1DD0ok+MWmAJ2SqwGBhOJ1RAkgWcOwxLBXWjk
hcQYbcL2QiQHEPLZsW/EQScOzndCsTdui8/qU2bhvWn+j+XWeHMf5kQSb0h86b3KqZSuOn9lpoch
qWV2d0dT0PN6m/wZH2fC0NeeGXbZtdeKDGQ6RA6vJn8RZuq4/d1HJOikveLkzrx3vPybXAPyX8PK
vpjoXBkQpylmCbxDOihnj07F8T2NHU7e6fl//nOCSiJ2kSgeyvctqUa1d78anpmYF0jHYwlZ74Fs
hQq+qwP04l/a5FKo1bI9LNsHd+W5VsDyr2ny68RGqpLoEQ3fJDtXg7GreHUjC9rhUP67mGYTMsbF
/UUsmMyB73X4KhSYGS8HCm8U7st5A+TsJ/LrCPWeKqyH5Wxdmf5FTwNS1M12qHvtwhmHp8lmwLY3
J4xo9sjyUQuglhMTROhynu4mg9cdu5IhMUboFG28LH6kiNoKraLWc2j4yzHXeQAEjI0kR7+T51M1
ppOBEt9YZkzxYdWcDSrkyqsxo3OdLD3VusT5/8tqDUTqS5DijpKI+IR5Nxg4/rIQpTMPMDKbdkkX
aB4pwWqaGTbC0+C1556sl8CLbMT40Z/xaWejtjO8uUngZQ2rXg/1UKWco71PM0wUwWzOv/aWLk3T
kVxII1Tgizne9ujw4UoXn4nu7W1wiO97DdUhkjJvi1io+VmZiRo0G7a6qxZWyknTLCpVHsAOx49p
rJ923kWY3X59VyEDSb/cesaX4CeedjZFpZELCK1mDrJr+SHuTF3+uHpmKALuRd9pRZDxcHaeuZ4H
x+OMUu1o6VItirjPlTkmYq6a+eichwd5OqHiu3kmnLP2CtT0F+DSmRnVP/1ekp9WnLnevbwce7At
dzfKxuDbk3g/E/RgMnw76o20lVN4QOgrdPXXHYdKjOcvHYJtfpw7b+nkUrtmkAzovwQOt+R2XmaZ
9pz9nsR2n0PFa9KQtvuuY6l9w8mcrjeqCIhPD817DDH91S1A5hFxoltVqNgQe1EBi63sJKj/sz9U
J+YVDDwRKAUIjad5KAkeUbU/HfKvrSsY6TkZLufSov284N3G5CsqgBjg4ixCKC5XBy5CiIJ0fZhf
sjPO2Fk9TkZudf+ELTdNjosXs6/riO3i6xQ+CW24eOloVHGVTE5Cgbwkwsp4gl90TycpqtTsfteC
XQ50ofmaV/dcOsULVgU/eeoUC7LIc+QQQfrhGTA0x+HtyBP3Rt2KvXKb00GkM7/X0LHZJzy6qlu3
ZU+s3VGM11uSUQJXGmlqs589wyCylQyxhmHXCzk6W1330s1hkREYf5DFJRn2CPkJYfKKOuZFKrks
mthVpExYcEDau1n5E2eIp7SL66eLNUd285q13SVjKnpgsqcQeWoGs5XjF4nQA/hJUYdH6Qm1vfQx
IqqVRJ+f9mVxyYJJ2exQb50+TQdopH0ZmCzCJv5QTwATY5NCMgDHAxNy6ls9zh/qx8rbfMT7Oc/z
I3nfMzz6AFs/XWQvA0iUYZSIs4G/PSAxMcK2/fNAtXsuPvFxBBhOO4HJhlwJLx6oWz19B4vWrkSm
3XePm1cmBeNAHm4IybxZDoGtCwYQRGwfuYfQlrT8x9RW1u1LqiQNOe4m0pYeNnwhvecoxOwkZGfQ
9dRLjvFgBhyhjc3jkxvlAQwzMtdlkrYIvpBZUq3Qsfz9f9FxWdMJq1IMxq2TFZCxOAWO8YDSabgS
nTyVB7Z5/2saj2F8pffczkUz0krD7Jx4XLQHxUqYSV19whLhbRqB79xYRy+uBWci2vdHqrcuXVQc
x97z/lNzdwKrpejnFqCqz/Fo7Bh+2NhVeUUbDSIDEPj9h6aTCjdiQNpx6a1vpXlhO5Bh0cKZbb9c
qsTRVHQEIeozUmYK9SXr5Wzok3Gcv0AO/sWWGXBxODNWqzUz5XLrcUJpBuivCOZJK5g2pLCQF3nM
CMVytvLFcvNinpkOEbp0SYasGSiD4thBk+VB+j+VkqwcCoCRL1/qfnnTptND9wHba4mbcFT1BfNM
YiEw00bkDwaFHmLXW1EwhI7qs4k7jNEoRvIVGwPh+w6RDvQKYtt5Lg3xDqB8VNeXfk7+CGGFsX/N
Cw+vZ5+exX2ikck+khWKhEE6cB+r84jWVVgFpDTEhBOMT6tRCMfLp+4vwzKI55JZpo8PpuUFSJMO
cR3uyETl0/jg5/LbOh5PiV7IpfFuP/RQw4ZK+fudXf6VPNL8k9O7S9VRwDTaOs8jtR2jJhQ8CQU7
jNcqS1yFm728HZTmkJok/B1Wtx087rT8FhW/EUZhkGvhQrYoWXOPNDqVxWMFWUAJiBPtwHFRKafr
dVeEYunUta5ex8caUUcTJgvJ7vL0wuFfo6EY8y5lYbUBbcDz1eYORAAAbx5JkYHbW2+VX0YsFpjN
b0yMznrPbnYMXUwExSdyyXwD36by3Hy22s7cf1mlrGzGIKSIEapSJQmBh2oDn5poEoqMNMbWl1bI
d7nsAx4TO1r2xikBe7uCHZXXR9EXk0rbTxfZYE73y4LxZ6dd3C6RjWL8zcBQSvvU094QOtIL95zD
DzTM7zm/VoRnx2hhkZhStQ2FxBN3m+ZxHqvqgv4vsGn4VdJYMu3dLfStnns0/b4aI+Pjrba+Q+iZ
KQ2atSmjlImLHNZB6DD8wGb3kXIxDOXfp+NyXywm1g6J4Mh8DN+kkWwEFp5Ry4Zl1LxyUPWnwA57
znnie0xHFH5ByrF+wmqlU2rCr0FlCR8Nuct0rq48dHX9ZnV6q57QZKVDSn4GDMOKD4BKojkLF+Ap
JLNYKO8miIqoc9jZBRUqTC9VClEf2q6ErJKSmCBrlyHBhNYzlpEycOKRVOyHljy6xEy9U80vvxSH
Eh2Un9/OaWsM4nV56A506YLbFsWpSN9dfzwLE/pkgfiyiFaIIFN2WL+q5A9nWBULEq8VIYeh4bgo
xwh335EuwLVu/TZe3hC2wI0sOWJSqEzhDyPNqj9ZN54bhDax1EniUEtiDn+E0MMMpeGJhj37c6ny
1D6oiU7p0m1NndEod3zm/+v3m34J6+eIEQmp0WvFtHvh0Y5ofC5Cv7JrlHhdPPlIn3F5HEci8S+V
iI2P3ibpF7r26u6UN3cIRm/uPWs+69nFR90kG5fphhYGcXY8/ZNRLsVAqrjtNPYzl7cD/HeskojE
rq24QNEy8PjMXOS4lI4JP7sTnNawB/v7RMNzYae+1g3cRqLx121UzCtVIvMg+nab4rmvBDg6hcjl
bSfW/ff2SWSUb1RsiL5UoZUfuAqZ5xpLTZSKSuUcChZBMwuEWd8P+vrk+AR0i0GFDXXrLH8HH/pd
wy0mGjOOE5VVFyQU4X57+jZaa72PadJC4vHwfCh0AQNOiy33XV+seAxSPZacrdnvGIUDhZgd0QAt
iBoaqVM6LzkSn49vCWFZOcOkM3isNX0yCWQyTailO3z+92yrBrXdkI4/cAIiQ2ykq9QWTM+XCAYa
Y3VctSFdrh5jo1y7u4uIcrwdcVhyJ9cGSyNy8QdwweL+AtzWFo2VMGJCUTNgpTY9w6y0hQmgkcUx
1C1hIsTJ7+kF5CfnO5GdrLCgZRJAzeXpNe20K8tDhDXIVuIi+zWw0hO5oeFWzfad2sIg1Y9ZKDUB
JQYrONn2fXgyGo4Wz4fJmyCcwTAxILB0laY9v5XpxFvRoLRXfdIK+9Ccb4+smtOXVfTUi1CnY0ZU
jIuHyDfsPkVWK2+O0WAFiPsHQXxhSVdydaVkK2/dI4P3HHZ6C0ai1aW2mT6D7oeV6mnYKFB3Ys52
cc4ufClkRavbuBTQHHrHLu8XLVZRdSyT7LhZs+TXg3g9hHwtMQy4RdWGsacfQeHVaxZwfchUW8UQ
y2+mItMoGXaS+pmb9gnaBpiK/b8Le8opzG9xBi1sUUCedRFLIsK7sErpM2qM6JARr2E3WXngejNr
sdC34+thNYRmRUafeKdEKckVUm8dFTqqugorK0GFnF2HUE6GujKwMGsiWW+0wpAMpICbNtdnpGt1
bfvjGynhuqkMNGvGR9GXBgcXvmsq1tK4JpdEl74AS7riYQvXcfiGsGN6y+jeMw5LtQppFnuODTk4
8jVBR4DnhsmuTqOoFYWuaxBkGTOkgnc6aiQdY/6ZO+niystK0jB+XnKDSoJq2B7FPQbbEWSLypxa
dLw0bI9qTN0pWalumfIiZXV0NJXObzy8sa9jIKIWZOftGWJjDd6GjU1tuHyte98eA9ut4gftNPT/
o+VX0fCj+6cQYggHQZEBRAGns8QP6/BbjbDT4T2oK9WQBkHWWPYW9OmDk0Y1UA39MeK0cKEo5tnO
NdkUAEZKoo0kZHOhCtEpJJwZKtII2pW4dYEZPZudw3E5RCZJ2h8fA8d4KeXQ2D3Yb0pODgosOxFi
fre03x/FDMImIQubppzC6lCAm/T8xnATvVPdVCrbve4YrPKDLcB1W7TdYAsjel0f1t4dM4MCCcQe
2ORPvp4SA4xi/WNoXsPhV+4vbe2WnPru5rXUCMe07BP06o1laveJ0nKIefTBsFZcEBmBpu0nyKr+
lAenm31J7y+wRbaXQr9fNOjnN8ffRT161zypWpyhrZSu3XA7tCDxdpRQ9aoWOUdsIhTGHO1PSW6O
72MYq69A6TokjiMMM/TkN+ymv+SgFjixDIl3wnYRhCPpx3i8tBMUNfrx0HrhQlq9gQnEF1CH2eKW
+OxNf6d1xt+a3tyA5d5x40admEtCRminvtuLIh1wBjsWg01FYz4tppVl++8xoPBITsXYTJj6M1Gd
oPcnD6IFtAYXARnCLZe3F42E4m7mEvgKyP/nSkoYTjs7NTYZBEY9RfPV9RgVnFVixizD9RU8b8MR
3ZtDv7Mf/QqTjZ7qHLbctVY6s/w7UNa3N1x6m/Lm5XbPAIq2jE5aagDeIiwRaCdGVcjpM3isknII
Ryn7MyX83BFvZAdkd45etV2NaFF6CG+dR0cpd/Kog8885w2hE0lhZITilXHtsz8PBfVXrJaWW6rd
wQ1aG9UC0Bt0vu6GjPO8/bLWAJA8TFWooiiGKDSGN0weHiJCtVwjrDuUbswTG1UZVtNBttGcp0M6
miNO49MLQwYZoM4b9KELStc0FoF7sQVIOeBQx87zXWy4rUxoE8c6l9hJq2KTCVpCN3RAPV/PUPQo
CYQazcLmeErx7hT1xXTiLmtb9wrXrHo/rJCS/ImD5wCUbqFjnXOi2iQ2k61+2xtepd/VCSmNsmDq
KzlMQcScuIVBioHJPp0NnG85oB2nWibq1N/WlDfbACAPy45enMGc0XaYNuD9S2d2t9yEvt0T+Ls4
9vUwhLnvCprK22qHySCVOwRZ0ikG8a8qMfV3mqnhRtXR3oVVYjhFSJfNWlVQBdGa2hF+xl8dCYDA
9hImEsXtq5xdrDx2GUSQ3V48aHNNFAdQ0kQKAqBMuNVXu38+A+O9W98w2zj2TUmywZpnZh1USZWn
i5KADLcZt1a0jXmGsqX/B1zXlnKAf3BYXMNTpI5wSQGuBC8rUDiDgOQYMRFWPQ5MjmQ5o5vmm4ic
/qe9AsOZq3vkIrRbEw78bYKXxMTztBzzCx2M9lf+v9oqpcXBki6EgB2ZDWsmMikkVOSkTryJdCfX
7pmYTp33jPzkg0peWSgU0nBZdEjEuPpLj3iJG08tUfwqKe9vgwGY7HvwIZ2Pyhq1AIf9MK+r0gyR
2Fjc7jsaFh9ZSdp/B12AKXBAXEA1kQjGT6aPcaMYi3dYZaCrHzZP+4qOIxUWO75rdnQWfRcKLxaV
TAR4EvQRl5gH7bedm3Juq7MLF/FFNTsYNWBVNcVX68g4QV3zfOJLWDydt6/bpgnv5Z5qJ2RtkAXz
3fEEVFdz8siA4BX4/oxWXCIeolEr0y7iRlwCrtoFu0o9rm4SdSOCwITgfwQxYg2nmHdkvm13IhN0
/39b5NjwwEsEPEgsSOK2FpquhfUi7bvtsp47XhTrIAhAWmH9JBi+eSiSbslNQLtH+Kb3toLW1YMl
Ati0Vg9NiIrIkL6bafxbUEyXWZUpGT+E8AdatZCbTiV+UyHBTkQ7d9T0kCOjPLSIeyGd0SnVtzMT
SSeY/EJ38uTKoVyEnPhvYpbS3fHeoYNisibQKqWIQbbF5d3yJ0qG9mL/FEJTjnXlOqTrH9x/cHFA
KdMPdIpY4j3iMODoozCrnyXapqshfkGZ0XIlUxhmR7uKmakgxpAA/Syt2CnsaupPrwW2YJTmKFYB
fVE8YmVbP6hEcutPz0QuW6llJMeirofYPSIhDx4Wj0ls+Tb+GtMqnTL+wzojkC8WN8Vv9CeLE419
Txxw2izFZV1guk1DOUmmOndskoxu5jboXqlZjDMeSDFkIILSZEZnza4rcZvaP/twWoYScUlt3Nom
Fbe08h4ZuCMiuHLEp2odS/nxnvmPI6XnEhCOAydNqr2LJIHEfgY3/ijvK1w7Mg4WsSkTqlNp08IF
PPGahgVsVNI0Pa3h2jldSsm38IqjpXGX8mZI0fK4DQ6pRZ/CrWiUxGwEqAUcAfrXderRQ7Y1xxYG
nhRSggJ+cMuuzHbzoDZCXyohQeOAUF7ByXPJQT7AZ7Nw32Tezdyewli96G4tr5n0vUcAsrjaoS3e
NBb+AGjmnohtQM2oi9TS4A3UJDT0BvjsCWmvS697P2koVkGAbphdEJcp3mVf137QGRIQxnmJ8ha3
tPSlps0+I6vWzWCm3ljaER7vj+cRtIwSyE8OwqIcu/pqRyH51MJrUqVLAZWSIuv44Ayua1eAZZyS
VES4jJHdMCSUlina8qYNsfI1Onarj3rVFBOjDtcp0MN1GdzaU1zPnVXFLNwuz5V1AGkIqct2u+QT
Q3XiHerralkXVOhXGZ8gZ1mE6fP2VXsdiU5EU/pijwqYdg4IUcJZY2KJzswKIfsIJtSt8ofvcIR+
Yd1JwHznVX/7NqBqzqB1I7ey9s1UalpuW1sgin8fHLUkxkzf4y1GKaDtywov4hIzScguKjtI+9pl
gYQa6OIF1swdic21pmKjJx/vu+mPAyM9QAMTwvZ0W48/tEJZ2WzOAy2vOPJJG9+XBSOv2hal/t3q
RCDqws1YS7+csMnBoM9kmkIlOD+KT+bD3fsgDwkEtLXJ9otkD0ykj9f8qoPtmMSo4mAhLl8Gab8w
jlUpmLsak0IIKWT4V6Z+bZMiQ5j1/tz+d/2TNdD8oRCzR+iUzWQiTr5+FLHqc9DAr7nz6uYaClFJ
s5Tmz8ba09VkGrxW93LW4zPScazSo3UDk7ewmGS5e1FQlJhoe3zBA6tG+gSO1x/F2GtcLJGF7N+M
H0H009lMuw7pZRXx1ErwuI63Kyad96RVdlvY5LKNdcV1KDcUf68i2dkApHIomjBzL0LBB/tXJ3Vk
77ygQkdAj5sY2Pb4wi4L1pHD7trS8Urky2kL2PU9cnBIvEo4Rb3EqKbuOuNPz0SwgWtYcSXRXS1P
XfTqZdusYnaN7o+dmRtBUYuSRfUld+KGkE8tYvfgZcnu02pc9jN0vUqAtRogyjVYLoBzEPs4EA6T
trW22ULuqh6QLSZeLhaAJ5+q2iAX3Q+xIjnP3W/xLXs6MihBYYQ2y6dgzSOghJhUSYjZzFn0XKKg
/4jZPRC+zWlbHGMqBya9LV1b/XuS6I3nN83L56FDBX5qOcCulUjgwWE/0olDemHk651EXtGfrL5N
UZb63qMxmFGkjd6aoCfaAC7J883+bOrrAi50UQs2s07w/GgzFQo5K4AqoqneZO9XvNIkLbqEBtAd
BUFCuSw4rqAvbjfwP3V0ck57OidatmEUpcrbQ6Bt/uHDQ3gC3tOPBBRU8FrHO602jqtgLXsDN5Rh
EjP3diXrVMWYXo2CEJ3OjlUgehA/LnhSEZuVNbln80ZOqfkzMtYtBO23sVo96lJxzN8NkEJBgIxm
L3mYxFd98fJb+KdEAYCcl0v2kbWqp/dkmtC3pfGrkvRMKcan1mAVrhRNfL5ebaMzH/l+qgxrnNZO
9CTdQd65VnZzIyaWj/ifto3nm67Ke+y9mWM1Fx4vBI5s7h/xwHC1OAMId2+ui9UzGsSAfqS1UJuO
w9nfVSYaxJmYXQHi5ei6ZgjrS6RSCHUSdRM82Vqs8T78Z/hbvrGv/2x8SlUEyzcoXv/OsR5rdMDV
JttjD8S58raWvqAUMrtS40P1wCa/vmyuDqTl5UlQ8OjwiDkBxa7x+VghbIM3wTddQngyaHLQAZle
wk0fXr4EYGk/WZarSDAlLfn4Zx71pQ9wKJcCrf48PW1PrtlJ0+WXe5lLX+trvViRK7QcT1QiAxpO
MVoeJfd3fy2GTsDjkg6xa0r1Oe6Rua/RDFaAs+UkLAPfRsetAGbY73gh6bE1Rem+e0dfQupHUy5n
p3Gnp+INOO40RjFTlF8MIfVCih6bzHyHrk7iXq19WQA8efB6faPDWZbDBU06+bJRpVNaFNpPf5gx
dJ/Z8g3wEUTWUzRt/1hq8LAQT3J/aWWiYKBYLax/3Rhf26wQuz3jB8TWzBMMDgUdmYQU0AYxpGDW
anbRrygWB0+9tl46jLLFPkHj8TtN4wk+Ak8ICU8sWSTTV7KeUUGIkAR6bUN/0l6EI6jn3UGd4G5/
Kp3Cy7NA1FKFLqng+tRX8kU2NFqmwFfSIujh62LD+TadU+7MWJb0/ENq2DfzlB7rgqljHMp49dEU
QGUkWPUGi/tTTX0Rvck18kP9zm9w7qX0G4xgK8K2FziIZ7brCx1m7uOAWD+P4KpD/qGvcu6cj2lu
0ooY8iCWyyEd9e0ibJvA/K7R0+IurM6Xw0J1+8zAQ7+NLlT2WPtZ93f85BVR33WuKmP9hIKNt6Cw
XniorFlzZbZtrDbctBmYk9v20/9cpnJRYr0AA+3Vdl4DPeaqdAMzNcuTOahw9vbd79cfBe7bIVgT
aLoDQ/2ctngsQJs5KNJRXoEXCQJzWMJTamydQChC7xIW29wdTbhBcgtCoS93rS/fJY00f38dcKmh
WI9Ef5OAA0X8dX5pMqAxl2rE0U50+5y0Fach1Lc0+k86d/7sR1MGgBPn8zi0FF9MvCHDASrcQwgX
U6MMJYnxXw1hgqa1iiygiCQAV4vptRPJKZTnaMgup+fAEsLYfK456mRJFGHd1tRTy78IKW0ZStmn
uBgkQ1Yib0JiEyzQEBYUKxfQeaLp1FM3YPUrjthzNXd6qhNnTGeW6/AVZ6dnM7pv3vdd6RZBBRqK
+6yNyuPz3SWoF6lAcu8ansjKlxiLAgRXIXD0Xvhmj3Q0R8obuiwDm1AfMnV7cw3HIepL3myi4o4V
UeNh5muxnsddMzoYuDSMCoxDMJTBYqQ3O1DQFap9WV0XghslxGgRp91u0FB6d8dub3w3OWmhJETX
k/T8nrOr+X7VMR0c66/fUhkLsDPsd83YcubMeVgeAzeinb0m68vC6ITVWh5oDIvNbDuPWpylZ+fd
x6bY9MNx8eVKwCFo3XQ+Qqx/Gjx76WgPb9b5Fjk1oMS1ATu+2ACXxjX+iaBcGp9tlDgCsRyPWp8w
wt6hXDAGoZtBNQWiBys07zP5ySuDQp+Q9Y5hq24DZvD7WabjKYRVhsATrC3/DdQZ6rdnMerHwW3I
yf0VPfNZp9P7XIxgxpLPPqPG4kROP3Qe8AB6SRowzwsLk2MT5rc/l2tk018Eu+MLtdIpFHrZZLfW
rtBPMxQSHfBnqkLXSno+Xy5xEb04ZQULL21ClebP5KNRM5o6yQGY10eH1Tr/IJks/BdaXqTD6QO8
vZ6jBTKXsBxj8OJ2bpB2QF/4A6un4dLHFwhvVu1SFstvrZKqBi4UTq0IEm2IlmJ1G1JiA89QG9Pl
TcodOTxlYiQHP6p4SfmZr+t8hbNVMTryzSjrKhaZQZpfSzkCgINE5c5s7dEl7cyuGb7kF6QVpM0I
hdYUaHU1AjC62blD7WCptfbvRlL9/dPoq0hdUW+xemH3u0CiWX2sZT7wIoQVAHllBrn/RRR6i3qu
M/7UmXIuUULZEbve0sjg5mE67HrsBZcyM8W2fzflyNIhx3ZkEy5AUIdqwbzdsbQEprYBSE5w447b
oCT9oLpmss+lKO+HLNLRR8cECYthBB1extjh9qOf2fOJaD59JoDZppBmytj+PtFLn8S4ry1aKnin
4bBO9/DgvtJ8A//8r2K5xrpd2VBbz+sMMUi7IwFTlJSmxIYCwprndlGOr6ZKd/bh/MnMm5Y7Jxm4
AMDXpUYikW9cGX4+Sb4BjLBfQ1wlUGvpb9ZJ6U4XordDPw9ph2HDfmn9IOdqNSUTK8KJ9FBajUsD
Va1QZW+b2taCCtNCyfRCnGGeslRG3RmArM+t2OBMPZlxkF8JmZVdGGPja+d7xd6/MVcnKUuNVL4O
TncYXcyE+p1FpUeC0plO9ZS3hxv2oTUKaoLRBZYFCNIjdi6srXcCNJQEu031eg01ID1gho0i4n86
RwkHIa4a2iapggkuutkwg1mV5GbrZh//o/Se9+Jgix56MGxsIGus9Pu/gvMzr95MFRlhpKwweH5g
4yFGfAgfJPacCcGHN7Bfp3isPPBLrMCFpQXs/AESeXl3PQ9VotZOWM6tImyF/8ris9X0Jc/kCGXF
2gJtfUkv1FLbQOa/k1IMHYJ/WMKqi1S4AzAvMtediw64r8p+9OPPFkRVRK6bevudCVFHaiQLAxvS
v43g0dwwIDzyWfuuqYj1+iAbU0QWsT5Tz/7xR/K8+2ZObhyHyR9vvVuGycZw76QSQcP7kJ4TNIf4
ZvWCOOK68Ukvy8epkg4hqJaFod9q8/DgKnhjBJX8YPEBguVgSTEvq1jiRNQlXfoJVE2/1XSwuqCW
qKMm5+IDstg5ofSxfLtj+rVP521q0cRqyf5ALd20dtetZvDFJf+BeOzH9Yp8kn72GRjht/zQcgij
h5NWUEHrI+JLf1uiBgvfTO0d+tcka/ZIVgpYVexbnbUytV1Hw19vXUBD5/n1d9dkn2Ng0LMlf2H3
NRX9sNrlGN4YyGLis5ZIEA+croYTP1CmmXKCtPoWARqVsw9fE4xfulfyDXbMC7owNK6ftoulexzB
JZP1xyRlg+ylXG2GG1tcZSRA4HY+6JND+vuXF3yksLK4cyOQJYN/6BC0GMQeApY2bF4jB80h5qfP
ME6B0TVIPAWQYZOQRwN6xjsFF1nRQ0skXZ0/dTYE2uRigh1PtGM1bTVxDQLi9cQb7jCBSCyL2ZPb
dy/3/0Ga/U6K1BoofqQ1bcUZIyOBvJzPox/6f2IZAsZ65uzVspKLm0QAfHRIR8dxQmdm5XoyNVCt
feV+rMix6FTEFRjC+acjuEl1neb+aUglzwNFhODOc0XVsJBNom6JtUBgLRj5Fg/87Cjab9uxCgjx
N49Zr/gPcGNDiq781tMRgkij75tqdMLITHmi9klx2uLweJdBld5vcjvgt63Tyy/E15XcMAzDxaMa
TA+gGvpSPhLp3vOz79S5z7j6kHz+CN0twfGowjbIRR0/W7hq1hQR6g/5wQkn2VXvBDkVTo14Iynv
23I6fDYzxnAqGeDJX9CE+lAPPWeJX5pJ3+z+i+EOHYENvo9x8XtPu+ggjom3uptRdF0uxbtuf2co
zuAVFt+MDNcSQHgXkxb9HEZaUrnxUUTOpF/rgA/FQbyaq+7/iS5muYyjVDQez6QqKX+4CDAOm6l1
IhNG2pJB2YVG2HtVBvy4zRIoie1WibwqiqwAeHgJ3xX7IEG1RD4zLv+fZl0LksR2D/joOSMed/CM
zMnaoQyhv/orsQ7N6EFKcyYys3TmiES1wDoOxHGFn+t1vplRMdpc/eO5RZfk97jl64zUYTxaxttc
zOFvbIu/f187vHLVKyE/CKBjhrGkZBBD0pMxlcNIUZWc7Y3nKnQ4qrd0sKeEHxoFWkfBIqkJzaNo
pDVKcqL9b9ol6LydgKLa6gHc6di3Ow==
`protect end_protected
