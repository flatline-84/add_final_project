// fftSpectrum_tb.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module fftSpectrum_tb (
	);

	wire    fftspectrum_inst_clk_bfm_clk_clk;     // fftSpectrum_inst_clk_bfm:clk -> [fftSpectrum_inst:clk, fftSpectrum_inst_rst_bfm:clk]
	wire    fftspectrum_inst_rst_bfm_reset_reset; // fftSpectrum_inst_rst_bfm:reset -> fftSpectrum_inst:reset_n

	fftSpectrum fftspectrum_inst (
		.clk          (fftspectrum_inst_clk_bfm_clk_clk),     //    clk.clk
		.reset_n      (fftspectrum_inst_rst_bfm_reset_reset), //    rst.reset_n
		.sink_valid   (),                                     //   sink.sink_valid
		.sink_ready   (),                                     //       .sink_ready
		.sink_error   (),                                     //       .sink_error
		.sink_sop     (),                                     //       .sink_sop
		.sink_eop     (),                                     //       .sink_eop
		.sink_real    (),                                     //       .sink_real
		.sink_imag    (),                                     //       .sink_imag
		.fftpts_in    (),                                     //       .fftpts_in
		.inverse      (),                                     //       .inverse
		.source_valid (),                                     // source.source_valid
		.source_ready (),                                     //       .source_ready
		.source_error (),                                     //       .source_error
		.source_sop   (),                                     //       .source_sop
		.source_eop   (),                                     //       .source_eop
		.source_real  (),                                     //       .source_real
		.source_imag  (),                                     //       .source_imag
		.fftpts_out   ()                                      //       .fftpts_out
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) fftspectrum_inst_clk_bfm (
		.clk (fftspectrum_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) fftspectrum_inst_rst_bfm (
		.reset (fftspectrum_inst_rst_bfm_reset_reset), // reset.reset_n
		.clk   (fftspectrum_inst_clk_bfm_clk_clk)      //   clk.clk
	);

endmodule
