// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Z9IrlXo04bSTMbzVCBjiHZyNyGJUektmhxpjb2HDbjHc+WCHvfU2EN7rnlIM3BZhT9nfDKd+poW4
k5IG0d6+rferL8S1o2uqfb+pH/cCcdB2ypzgIh7sHa4FTmY50Q7QhOb+LUrZNG5AVk7TbSwbTJhl
iigWZKXudwwkcim6gFyG017qxqhp2WjhVFlyH3XYFEksdhQ17YIM7sGyNYQub2FKuBY7kDU1n3lm
HsdFyLEF2mGCR40kXCts6oDrXmGGDVsj/aWkcardagPZSHYqenYcuZT+ZFP1azcm3DxZCP69WLEo
i9jQe7prMBh6Ah5vNGeoYc6kdo8foT2U2rionw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11120)
3wvmilDmlswbbevDA4uCd9jqUmaIqrpH8y0QHuWK1B3n8oVA11SKQMZXbH/o5PR+OOSxMcLqsVY8
xWqTdPT+q8KSFfgxXAaLHByidVPwji021RKOSv36tcQchuXHOjFhP9HC0nRUlTDrhgCbG9H+WFj+
Igi1F3lwW3rlayy2/gTGxIXDZWXTHYNtB4rb2gVhg+43UYyLMlCI0sv8XkqdQIJdx9/w1uMXMT56
Oj5+Ojpd0ls2CHA3+onHnT19v4PqpaxmgTEXmhYeiQZRT8E/W8U+E2MNKXCWaPeZfVC9Tfyt/AuO
t53Y6Gu2Bvx84H3ag9YYTSc2gilozcLYh2BsVk1iNHHzh9pMD9i5zTeVVLY1vQ5MrXhFwucGSpb3
ew3nhALv9+mT+oaIJfK6YFoVNl+/g4KUSkq1aIvXFpaXIr8HA1rvqEy+iSljP4zoiGVLxo5jvuP7
xH2FctXqEJYXOCp8km4TFmnZlNq4nbPgVnrxSJ9Vi8NGN9u2VvGLLs3LqlKxweGVTnTZW29kRqLZ
B95WvZYLuG96X3M0A3IXxjT7hZggBFikXyWf5RcQS4VQfDfXk1ofwANBDpNZmMBF0+Yaq6t+uHcs
IuaB2RNM0LhVtQJSrWfj3vXtehJm/e9xGxfNIrm3MF0KtzUjduR24hkQCelm/gqflzHz2Cwh1z+M
Iq7t8TJSuGZflpxzCUbhWkODX+fLloORP0Rv0welgwT7WOTVIF32aJA/0CASC90e2qHy+j6c6Rfy
cfDsDVpQSOWetSCtzebXZW8z+PsxqWfIUkaDP9v2UXDJCD6XExc/oIkWjkiuuBoaFt02Krj2J22k
Tilxoiy7mx14o+Y5ywCJPbLaJCsYu/hkoEBYTmZOPXA+AdOMgeZ6E44/8Dp4zZz4Qwyt577vO7iS
bg9OIKjTt479VyP4kdqaKWieKb379EvfmKWT+BSLECsVt7LjPdfHkmB3c3nz0PeEW/rGeNriQd+Q
v7WCm2MUpFXVHoa7KTgpIIjGeq9m8TnADln5J4NRHIAcIaJQLMAlVfWFHd5CgIAwNucscs4felrK
03heFMkaoXuXov07W8LzIv5rtWI7el6UtX4rv50HznMxNnT1/0kWqVgmc0DsQIx/CP3dkkQxws+5
M8n/86+QgY1inH/9HUbdkFeXkFwFeg998z057tmPEq1TaXDUvExaDd4XQu0c9zeogwsFjxcqg1VU
4Qeapsezu/nJEdYYv5s4YOCpB1WidgovG16bMeLBKQtCyVf9FLGMYLoAZdVuEEFQahI7qOVdmldy
QXmaPhJgzCifs+yVpqvniQ/aFVVapxz9CvLzS3VCTX9mEY1IF+nayUyFz2diO7d0QjvNUHp4N8dP
tQg4VzUxv9Ug1vf5FjEOt2FqvGQzh147tKidGcDxw6XyxAt3Bvja61SOA+wDI2JbyONddMMZXcis
QAJuU1v0845Jt3tuMG42zOAbycWEL8ojLpU13qGApNPtUji2tcM/yC4ayslw46R+/nCWym/VtaA9
qxYgdMeuG744zDnRnxIIkTYLZD6ITzkz4EsYHAcmbEamf2zVUjQ0Je+nZ9g4Vedn9eRP8mfgTncG
h1ko9LV8+R1143yt5U5Gxnkpr+TerAChN5scNC93vHErAjA4NYx52/yCdITAr2ucyrd3XuZ8JVDE
POrTsG27hXUcc8HFIqMPXOrZUXogJWRsM7PqFCUSu6XQ/DOUBOAGs0H3rW7u4BJ0MrBqI275R82G
5m5HBx66On2LxURIpE0wKIY/3fLVcKyrYkr9LL4uuYi0ICPT/KuMbj+B5IUqZR+YshDo/VtjsRtA
Uuq+lrNNvvWp+3/K+qoAvi3wVH6GKKoAzmK7pE5wpGe09QfD5/5LRko6ZfjUqFkFXaNyV7DRKWDH
dnw1Sjg0NcQS7B1M+GUys1mabwAccERRr17u666kd567gEQV7WmuG+Af/KbbeWdHt3ODDl65tzF+
p5HM7uE8plcMk/ghfbcwbM7DNyuKhNQF+oLODw0afDh9cU11TviKmdfp2irPOBVUT4lV91hbCfwQ
O+IEWGewL8gFUywap7lusNXJeaRhgJxinxS+KaImGnsX1o4Bm5cxxpsYwZU9rIabVY0lFX5Rn6u4
hEOClu7HSljVOqRIIjnEtnxQuaKCKcU3jUOCDyMkg58MnqBaU56o6CTP6k2kSxGznEkMIqurW9uB
EIHssaX0CfKfdg2dqNY3XeN2Bg0crNcgXbyHPdIlPTeG3bFEZvPF4g1YM3uKkdv46BVsRGutDYyz
a5cuzz0fFLx0ZwBxogROtxYPRRG7NyiHKpAH9hABrIMFh+CNqQYg8PrQQU625CW0TVq3J/LTpCuY
IbwyTnyui3GKTSugsIb2kU7ycAgOSU8pRD5iHIx+EE/yB3kcoDW1rLIdaTLbr0Bz7X0+m4gkNvrR
C64qkR+BR7MV9xQIab1/1ZS7QDe0EKDl1Hn1vt6n7H1xdIfLL2l4rnZrbTirRc2nzdC5pZjcd2wq
20/FPVOk3Ib3euiTuwruFGvQbjLn28aWYDGGecZWwQGwBLJ4cSkKgO2btDlWkF9DBwk0yG0jYCQF
QEFdS9nySdi42Q8shi/vCOfzK0qqjzmfuWYF3LPEFrwcaQP8zk0Fr5rmi9Nc2XsdcgknB5Qxqn0d
/GAjiCf5wNt5/tCbpkGKmEW0/t//vTxFzHswI/deTSSefcQo8CkXmFGxtZyTPilQOpPFi+/oYhFI
vgXPJN3WF0F8Beg6lsP7DpbdwdrS78RkLS9l9c/JakjAaGyCRoZmSI5FUeauCriN7Xbk7HtEvmEL
wbtmgLqzFjwSryY6eHnuZ8WqzC0i4ARe/W6s9SUYEaEu0OGgsuo0u2pIEPKB0DLEMUQCNKlYQxbN
kG4KIWut1c0lFvTk7hVEQrU+zhxMUxkOsgqar2LIJpaIymalrXzjolt8wpHGHCpLtE05VxnH1cXq
BNoLenRq2KSUllJJpzdMLUfAORBtNfmiZulL/zY3QzV6rutOo2XlFh2J+wpoUR+6SEjnZFtuZmy/
XLUQOcfY7LKBltKZyf9St915tmgh5Ncy0Y/uhZi47/STSqk+AiSPNs8suGRZXRu5aiOgB/klJ7vL
WLkamJ2pOPiv2aAlDHETv36XI4YUV1irpLl2VkZCBNq9JWfZigG+RPia2Z0ldJChocSagIMlBQnZ
++OYD6rraU1TbAhVqrRcdudlCaMdeNWK8T23axmNRtn/WVx0drdnsBTYxiaOIyaimMmhUAG+b4VL
MFwNFIo4MX7RL2wSfb49eYZ5B4N+QI6141SjJGHaPLJL2DBR41EC69ydi/+IF3IiYMn7gtPZBK4I
r7zzdU9VwGTaMuMUFC1Cgf3te5YN58C3TcGuzh3vPm7Ig7Ob2ZVf7Bj5POH4pD0kekMn4XQvOGDC
L4638FkqhSUerYWHkGS/3WLMjh4SBYXE+ImBa8T2yz7vAK52i0ZBY6x/2kGNumCAc6R87LE5tCYE
qqSAkCHqNWcgb/ZhmaAdssyp+mGfVwe1tVSkfy6WBK9lNL1ia+xULZZ5nwFPb1dtdWHXGUN9ZO/e
3jTM/htbdRB6oag26GEm/evDqz4SjHDp11PUbUSIZjzbfngMww8mg+jwN//vhdkpBrUKTHFHiG2I
VMxOfUQu1y75wX0pUIegJ7KPPlXqC0nYv6xlEExXg5RvH8DsYf10/FLa3f43+zWXrAv/LgoIPwVW
SWvYzOUnCqA3ARo6zurVfb4L7dv9pUxvGYLiI5lQdtxGLpnVtbaXy73wm2ZUurL9Ms7KCW5SQoIs
8c61w3OvQksDXyPlh+uTI/7gmumBEjZp98wuZ3vvRiilKsB89nSPrAo0XlhZpq/jixz1htZTL2Wm
SZ+VvmFJ7UJr8i+sMDy0T6HPxFRK8VtGd9EVWemc4lSoFPvIwm3xnRJAZIbDB7HwjSVLHQeTGL/Q
hp4GZRw0iu0HHbb0+akF438mXJwe8g3aBB7SP/CyKDJcN0WKyyk/l+s9wFJoMmmWcoEVO7zCfNwo
Vfyj4hVAE5RHj/mfXbAvxVY4CCQcZjg7cmPCocHoQNAY5jWBPKPbJk7U/GnX5VH2zp4wc3Wrf6BK
pqtj+RPM1pn135bbaa7A2jMwCtcfoz5jb2cLpGZ54HsdHQWZxa7hK02qAlut4kRL7GBACW6ql3yX
gcgf1cMvy9Po6VqPeJr/IGpFgMmS7NZxFkFfdLU+QBbpYWaeT1nrwYIWlBhWKdLbOmPo/XDomQ2t
ybZYgb9HBnBTvXyN59E4FIB/CYpw9MbPTy5InhVNd77ksICIjhwFFSG1pIwG7ndSYjcjlok5rGut
RXukb8yjExz2rSHsy4JaXlD9Kni+EIRVfgQIFU/O6Meinnr4h20B9SwGuBpKGMFoBldwnOq/6N4s
2GKiYB31FTnpwGcxyEhs9Uifl9iCgIZ60i7IJxzF3RROlfOQ9Q9XkSlwuDZR8UDXk8vex3/Mbkw6
r5RRYeMMiEba8rjkNrV3aml//RagYEqNMTdXguvjNAX7H/t0IrbQywTcQfDV7+dEjtnvTkDNpvPx
FvRgDPorYHCzY1CkEJc4Lalzn589oZlC1fdibH25MFqcAPF7kX7KQvEBITihyTb6hshWBQV4y7/7
jwrBtBKF3puodALiZMRLJK0JJimSB+K8qdCj3rNFNpgSKgy8H1Oy0Nkla878Hxz00eASnXjeQfMM
eyWRfsm2Apno4i7JpQwjc+7zad7g4VTfHQ9VCLUu/CBTPFhEvcKjeG1I0gTakcc/xoFq4W1QaWdq
kXHXdEbT5LernicuWXiJwH4eCrX26INOHhMAPca1+nLdGSC+zLbHPbD5xykUQ3MLdiImYr+FSm8X
7T8x3fQUFUv/1W9v5I+SnrK1Gmp42gg1Da8bZCjGQobrUp1Dk8Bs6V6mzFVpEhPNoSsWDCxZ4BvU
AKx+TAR8exUUnUAQZxuNZ9CY/fhVknsr9r5VWnWDOYnbag10SYt7VVVvm6JmG7GJVStlukNth14p
l3Kl8Qhro5XaWHFBDrv07tRicVIWAXgMZp10Wsx4Mj9t1/avjraeZuqu+2FXw00YF1gKaunJU/Of
hF5aWMOZCbiptZFqnu3g1hVX5GyAJn36c7GFOhrOtQSgz70X2PjdmA+IEDSh7fNGlKmxBo8QLayg
Ui5vBY4+L36aIXXpLJlsBx5GiFCvcd6TNrLF1z+miHbxdq8J0sL5Yce43GiFmYnpDUR0xkkxSqIZ
4i9OtcsOvOLx55GN8dL+G6z60uUF1sWCZ56JtH72oiKJ+DB9L+1bs2xQDeJ8+xUYGf3/HpCtWIjG
vKPRVL3tmCSXYTwpPmZCbEBmSnK+e2EcmWcypIP05ZKxNmFsttqww+F6i3U0hYKrGXlXuloY+ntv
NdOgcG9olOXqrxY5fwI0Pj9p2VWu5O7euA9BvCuHAEDT0+MSeWNpgF3cWJnBpqx1F+4u7aILBeRO
v7IyTdaOn8C/LVDOt6gRGwF2GK2CayFY8D4IorRMEA8TdY7x/JPo+ZMzdlM/xwVTD2yQLWlGjSkY
tN07iNqFIpRw3jghTKKi3XLZmKEKqanwQcMEEK8L/TK5UlKNjDoXG8mRCfR5OxxcvqYd0gQCz8Me
IyCYypUX9YEIfl6YBqZcN+y+FFywomWpRKBlNmZIRM9eA2BFQcvvjy8DtRztoOgLdvqFLQVOjbqB
qxLKw1C8hZ3c1nbA2IJzvDgObH3yzTyhSH9W3VZ9lylwLVFTr01cjgOawTSbNbPfcD0+cu84sZWx
1zZh9b9+bYPWLMzlOSQUp6Zy7UaAnI9b3bsgL7lPdV+mpJ2NWAh5jtOcixLU39meaQJBrZF/m8bg
fmfoexpKlshC/zUj1pLw3nFMivQDQDcIecvqBmNWSvifPiPx2A+oEKDi/mmjT7oS/plty8NcH+Bl
lIwfFkRWb3aFz95yZiO/unf8yHknoOuRhPOstk+lzqMsya8BmNFSp16Ez7VIqYXR69h2MxV050Ae
Sd751YzLoRI9v8hduNcBk9SALZWOzspP8ugQjR4W8bcM2HXJndHGzl9WGyUJk7AQYinMGKbph+RQ
kv/Od+J04zMgJCqXCl0BAvWRKuPXycpKqNL1Yr/ukUSdEYeNEIcSQBPXglIZlwY8ix1RA64X3DNh
a/eQv85KiZj4kgtdQd0mg5BS2u6Laal9jLzKo4mLW0aZp/L82lzzv5E1loeobK4rXJM/6o2VxwPo
29O0I80bTH7E6ZAZH7ssn2XWUS4AxV9QM8sRSDbPPvECgX5YPWr/Ha9CFirH5eJqjVwfEO55WGwE
yIG2GTvpl2lCmE+Vnqrhd5fpMhQWbkzhfnqMmsQQLIy+wdAIkXwvNSKs8nB64Cc3x8WJpMrcg+W2
wdiscAQkIJ7h2atMagN3NoJj6HeI8xqs0XKwR7rFDxMSez9N3ecTBFFC8c6Snojs3Zca9gyJ6HoS
+uigeHejpHrp9bWlPK6P5Kk64KVCEC/EI2YHaDbGFF41dEanDhogEicDTiJA8+LNLiL8FlXy/uVR
rXFLQrJbsUsTyWE+690VFo4G8o/oVVGr/8Av4yIZi0NUIKusG8pOTTvnbXchAnNKe5gePEje1e2N
RfbdH1E0YfBF+hE1sKun93T/uA6yYS0nQO/5zEMBix67dB1eMe8p08gROKUFvoCbCavMKJGKscSj
o8RpiS3FXZSqLvpqdzlmzP0t+r3v8fIzzd/Ayj2UdPZ8HBDCKmprzYMH7kgLePyTqttSEzKlJ7HZ
JS909i35ZCPB3xYrwQtDSK7BUdVzZ6fMo0ktN17uBqNKG+H0kWV0sHmTXQVZjD3QGqNytxK18fJ7
/3A1VFbU11oUgpEMpBwZAMuAbpBKpRzXhSOQt8CU0ZHvfRRQ5Py48JkJS9+8mUvBKOoLa2ZYyzR+
wDdKmo2Fvd1S/SWF4os0jhGg7pxKAYJGoODiIyfccwb+eeDidZoamUDiCppIMe+2n+/a2ULCweZ7
SPCcI0nZIz0E64aNeh+cAtBnz4qe5/nDvwLU4YF9oGt36p2h6BZKhSfHUglQB7ng6r6v9xEe/Wfw
XaCmthV/QgySPGGCDB6eY6UzVGFX6ohkTR9JlVlsSmOGRTchIBnBAsD2DYRzm8ONylSKDYKC9rVx
5akdCzWZNyUJ0nqB3q/8ENYDLG4DuxTPJWODXCeRldjznAhWlf5UQmR5DBboqw3dgp+rhyl3FBh8
vleeCulQjwyTLEkdLUO1QYb2lD7lPIg3bVPdoQSP3Lo5pBtrE3rK3m9H0k80a7F9eMmXYGuhkmy6
I99sgC2YawoIx5MOs8lrBZ0xEaWHXSdY9/L0ydfVoRP1aRX3edBcxIhO3K7EuZn/mz45j+ksSyNB
C1COTeScMkpn6JUJ53kp5twUOXmtkAL6Ke4iEJQRb9wkYqF5KZ+aERJiiuQsnYOCvSCRUB9IpwEG
+b8GHrX4WFuoP7sg8AeJVHA8yDSuTjbeqURxP2cyT04DDAd9rUUoxutfmw6MSUhWwpLSHCb2ZJWc
PWYCdHYTkDjGzqsFHNXaVAvDczWjfixHK9cVhWtL+Xqx2oc3A4iu1cb/A8DFcCmj6lgX1QHFsghH
3kyrCo1bWNK8iK+w+Kw/SDXdHEVDaY+2vXI+YYwqVcqUHURUX8I0FlOYdndSGNZ3v0ebwDXZmIEb
kMLyJLQcD//50DmU9cbGTXC2lBW1LvFPmw20tI4zBfm7ez/k5wPO0Lo5W4A+jcqSbmXhLqPjqVgn
ngzP5ElJIfQFKD3VULdgjqNtXXT6K0r0roRMWKc1Y23l5s3CEqquhg7xGChw4lks6zsansdofZE9
YRyyR+kyO7X6Iv3orMsBkQZMq0Ewwjy843vYP3ncRnBrrNdYkXDyprKzARPB95erlMsEU4ebNDTB
KBOyhMwWhnHfoVeek3c0UaxuWMbNKZEf+n+xXrwvNsYrAZmKP9mh3RqDkn8tWugFxdgCrWaD5f8s
w9Oa18ENtnP6lnbvj8cs5NX9j4OciBDiYVNUG/TwCKxDsB8CbL9yanGhdAgrikkqdw7BBYcVgSx0
CfsffxHRqVMovPLPyTwhFFCWIjX1yqYPceU1wiRJdtUsJHiFY89C0aKN13UPLrl+bWNTGcsKk9KW
sRkKYTEabeqvtU5D4pgHhwbzfXfsv2J5UIqTOx4/iSWQ5EWQgiJ7qMcf6VPU2bKlb+9QUL7knE+b
iQgi8SiFg9dU9iZ2sGSq/t7tIswxxXjvAkabj+OaFzv5k5AOy959Dczm8i903rfffbEzB45+xkFB
K5fP+z8Spt2DyCr777vKDLVP/dcDTzmh4/UqssCYXlQBnNbQ8KBOSMOYoZXvnkek4r1xugMcnIbR
R1D2+ou6DTrdIRNIrkQlDOCKg20XypTvI9pTnq5zZK2kPwiJMq6gT+W+obaAshWuci+P7zuDpxto
hb2kpoMQF84c7ynuxPWXBi2hdBwenzgGiVJbyNhjQM+Q3697de9zj6F3toGMCANEs/LeEkruZP/1
sF/xiW3BOfauSdxjRuMAEd7jt1o6LioDIgRcAkAtkH/U2SCAz1L+zu9+hCL7J+2PFJBdTyYLsz6/
S/pPZZMSovHpc6XT1lRXRSX0HG+/eZHZIfr3s3//qDOAU03daetg54EMS+XF06LVkxS7lELK+zIc
1cnXlFiiJdh1Jphx56CPSmsqhk7q9Uv2df7Zpx3nmjy41yPQB9lPnrd42NpX+EPhfnD9+Jsw6Bip
Xj89dT2fHZsM+XRnB1yZgswO3fIqS5CSmu60eGzUrM6xt9+n+ilvkycqALH+mRA3Dv3kOXCz4AUg
iMVzVSrI8zjzfR80m6vGraTJQJOb/TINZXudebWQc7C41QuG0VLQ3c/Q0KWnCpM3gGn2303rMGbw
Q48aH2uhosAWEg1asMQHymmSJM0/j4e+Y3wY7C/8DJS1aoCr8NyxbPmlVTuKVLfzVkNEDtLRSS2b
onj/9BCxGpLrdPcT/tajjjNrU4/RMTBuCTc175M8gNTEN3o1Hpv63RUfkL8BsUa60jb9vXEgiX89
bXrLfEbbbIO/B9fPvl0S4Sg+i1+OxAWjMbK5wTDbxschBjD0MEZsS8h1bbGF+m3RcbqmbV1bciYL
X4MGNjeZLN4CVOIMMxaoTphFAYfYLE6b9+9QaxB7Y5JOqIMr1D+PLu+jjdncbZ71JMbJCkX+CUkN
P6lN8pAauPpUxE21usWGY/IRBhPyitS/euFVd+oRUYoXcgAm2tva9MvHCUuRG6CSW9LMaUo0b8Oq
W1FFD+Vz1FuYGo4CJ5eG+7RbHJQJzcuOIJoB5Rdz2O+56lUwwNF0twnI4Xjhy94ASJ1Wo6MrRjJ8
swgGbGMXqpM1wE4Gv9euMPLoYnJArdibqRrk3k8LGLptknGG66TJxLEdbrR2XNC4EuHSwDwBqdPC
Xkx0ZAV+WbdFCLonfPdqBy3q1Pds8tYK4QFXWnm++OUCfm/sM4RX+tLCzWeCJscS/2hymvXkEib7
c5KuAi0FPGPAsjR8JnPMYOaE0Y6haAca8odPEDg2HdNGRNlBSfv6ifgFaJp73RcDmGodahmMR0Uq
kkHTraWa8GweTYbJZWy2iFmGC6yZQ1KVlnWfwu5XyWSjPsiJlMhRz9I/bvO0f9SIoz4ZCtSl68+X
IQaUppHXlCRMrn5os/X91y+5/yCCxGVDC4WUK4Q8f1ZucfkYl6KyJ6Xn7XZ9zpRX9UAZaEQVL3cV
rQ6NshxhN5u5oKoyB3u9+3Hf6B4Ap65mKkSEs8QACeapEG4XEQ2x3hZtWviVaK3Y0H+2Qvaj2rVC
RMti0NanREQOxOjgTYMk1eJ/+XRmMSg1C06DX4Fq0KvC3CILRCh2laThUKK8STGWyeE3JzkECgNY
NHdxq86V1RfRWtBmy1GURbYpuyQqJes58sZCQZhhyPtczhhmaNm1IQgpWVbdDrtaevbCsgUL7sLd
WCusvODimmyOcDi9RO/2INhI1tsGeUZImBEmUG1orppbUmqfxhYmtRM4Vrl1ee6F5EC/zSJfphGg
CIP6or5GqsGt4KcDEYoRmrdtlBBHNjR6E7YN9xdqH6KQ++B0x+3+Q/wBY0ue6LIJVJCy1YS8COJ5
WkZRI2h0DkuiM2m3LK46Z/OOl4F92EZPQJDMlgPpGYSKlCahgA3fUJbd6eZcAnuEkaFSbwjyvY/1
EyWGyQbjyavGC2a0zk/xZ38hOTrEyhZUP/0cTpn6pU/CunM372cd0FvY8crgjQEFHfaxharKZK/W
/XFggap8eLvXAHtbPsd5BWgqfHTrpIldQoM2vI5Uamb6h9H2pI6VWlcfJjpS0/ktLgxLy4zMzq1F
69Tq6IqdQb6d9zNL9wpbEsSj6MFtoDHQEYmASMhYD/vqrPkfKEO6IQoDsdzmsLkZQ3nOjX3XODV/
vcpLVP9h63ALpvVj5oML/MKOYslHkYwsq8qWQ6RYuQJieDnKFz5si6yFEzJdBGJfTtLgqIzJi6CE
lieQmuVo/6V+hhTzSXk7QpEb2+7N3mss5bNycG7/p3Mvkhff6vsbLBm4nw37zpt1Yp5ugHcK+8GS
krcpe9mjHpbKtuhw2U+DlqU4Q6UUXrMZE7RkV9KcoCmXNoqRSC4ITsLvQGQdRVYLA0EceKMygmM7
/qjCgROOuzTCnaJKNd37EVXrv7fpfkngVGY6H8RNEBzBYIPYzA0DL1ZxloKDI4+rF3cRMhGupq5d
pfkeccG2mddtmcwZq4tCsuoChOnUzuGBUvzW8COqq3iwP3/z8k3Rbx2QGC5mWu1qoqi74ChBLFOf
zML+HOkJaQIs/4nsyn+AyOOZpSml0xBY1Jx7H4g3i2AVUAcgwCF6juoCqNPgcYlJrRr1RynxtIck
yo956eYarmZXEMq11TQUWPM1NS+yLfRALT53UXun58cDddTopo5/3Uo35b5+/0Y3qJFOD/yhTrV4
ULhv0SmuOMd+WbwSwuLCIuQmPohTGOuzof3JHtnOnr4XAHfdQe16qHAY+Xu/edcV4uJLndvhYFi+
XKPZRcrFtkTiQIQw5npdEJ7ejXJU3FukIfm6n4ftQTlfWZKr1wQUpWtd98Zv6xBnxnjiDwWeJ8Le
Rq+QVREPQ+AlgRPvH8rlVbqSmcbpMn1ROtSouoHajsJ4P7w6MbuHtMZ+Ni+sCp/LBcrX58VENbbu
2LlCD/WsKonUeOx6dHq2UdVWPTDZt3/X67WjuAeCJT8ELCpoygmaP/tulSI/hSoaega+4JQor0Op
XSivAMgUUCKP6k/FA33O4Fez08x84Vw7Ybh5wpmnmxnU0acXRkkbkRGCuDVfKXEWEjxKL/StTPyn
b9QCVJUOvgjMWta5dCX5NlbzWraTsSpxsIQfIeDSrf5RkQD9T9L881PSK3wLmpUy9PG7xMsskjsz
sMqtpmyQaE5OgRGzjssZ+3FxpvBI8f+9mOsSbuYlIfYw8Cpsa/nB8ae1kFuFJBpRa8b1UPfVBT1B
99yQwh8VP4SvFKD3TAyVnhjXndFJcMBba1RqNZ+RdbkBaVAkdo96VjwoR/NRit00K2sD05AxHI3w
EbcByQmzczpbt9wf4c7kFSvDCPq5Yi/ZF9htFV5ckxXk/zEmeFOmO0rQq85/485cXp0JXI6vAGvW
Ss/qAHPuNIMbpHoFCgorLisszCGbYuYz8qBVL+bZJTJvvqNdH6zs5Cqs9sgYvkuIRNnwVOK7o02P
t5iJRXAPP99kiXVy7kFymkVGrzGjgqP9nSZbV3bsiwwY6oO0vLPgHJOlCv3QdbNNHmk+fFRfs6rj
fDzCTPY0WWKshHkxv8whBkZ4CN4SjV2xXE/F5SgDjbNbIydojGvrxfn0SpObRVh5sBatyZJee4nl
MzlNkFHSjgvt9PYZDPp+jB7tEa1x29DaiT+82+TBft9+jjTxG1uQxnuuYDV8khRHtyCVpr5JKqfS
8wMdOdiJBrydp3noAotj4qPBJjvQKjrIXZvaHo1ZEU+4Gv0K8deKggj00J0X54+P4HnH9XouvgOn
QfTgAUWhfsbQQvVwDPWaziI9oOC+0TaPmZ7UrI5A+stVWVz5vi3KZrc7hhKaacHdx4ryb1lVfT+e
232l+zqCFvvtDnpNUqK5SqbpfBNDTAQyo45z4i0tPWWXr1cRGfbr58C36N3/DUKjXNb10bLqYE6w
A4FWkiQ/gJttGaIjrxfhPJalrj6Q3QOGUEqAgQbFw36Gku4OeMeH2lNC7HDGdD/CEcMEGXKGcUOQ
EHb8lLlvK9Vg5ONBcPiv0gF/XFjyBbcFb91NRyNcXNds55g22GInh+SpZdg4QQb582KLhGUI1s33
oGLTXtjpwndIWrtWJQWjTuzc9l3KgXDKpBlKGdiY1XcPiEj/sxv5Z0RlVp4h1nVPbItcsQ5dYVHV
94egli0vr3USNP7pSIqlaYi/wiTAnQTLjgSMj1s29nfIxd2UfNUJo8MWD3xcFRLIISO7JkYrHToq
3jlzRJPAnkW7YLVvANslmVwmF5NmztAvzpGOOOV+pGoj5Kbvj4jU8JgNGy2AW8EFBPtWKI6+lro7
Ms7gfwm3BCm/P/oATtae+6+OQY+RwYmaVlbA25pzvoAxIU+n7suSmWmGg0FOxKcSfsnT4zRT6gVj
ttuvb6OtVjmFOOreDNPLney2N/uYdJ9JzDsKg6jfpsp3kgWclvfjisA9wazznXznOq7KCyzXs0vx
6p+Sx1W5dixQihtxJty2sdA3GwoviNLeNeQ92oqO6Q3hAA8fLj37MTtnb6xwoPxZPJgk39OBbqD8
elzyUYLePBrjO9CAvWwhW/ZvLL2Of9slnQ8g3l3Q6KuOutKqOqXksAfmmLQgEcV/cjhObhrpSFtz
w/w5rvcUwg45iAYcDkQON65oj2Y93oZlO2h3wnYVznEOfvb7yJVZufH7z3nMqCrPHhGBBESHWCBs
5mfW51NDpi2FioFEDNTmfj5MzgyvQodk6DfTB+mjQyaKkCot1YijUAqauwwEyuSFKcV2aogHMDg5
aVfF3kPxpzuR2c+9WpXRWIGuvGDVbSpNgkY56XkehxGc3qDBfKiR154YS9ILzzhw2w5ev/Nra41K
NjsQBtk3ojD3+T5eA8YHB0KIft2nb5IMBPM+UzHp8uh07dStB2Wq8cd4DrbOHwqJUY7LzdMw79bT
Lc8eORfuPwkT/wtiwTISDi01UJQfkQMnM+rg+r4K+E7JdVkoP6cMHi4e1A3v8rxr+mslA236StKA
xely/Tjo77S9CwYhS2RpbxVnsW3vYa7up19uidt9ubAp3qNSxNyMoJMprH/+YouvW3PvYNcvZKa5
K6AdR4IIUcZv3vRBDFqAnanZIYO+ID27mLZsE85IS0mm19rYcn/ZYKbFkEhugOb+aExAIojZ6Pgm
zSEdT2GLEJM8EqUpqFNtges+Mpl8fuDDgqiV0UsPIECPsPYksnBII0XoA2j4fr+CuNR56VpHTHqm
Ad8FDVztL7N3argwnZ0m6HYxcKivGs7eRZEf+fGIj/5BnUvx1BBGauw2vSWDYFIclSZ00dzSKb8D
XMxZ/LhE849+JaJ3LT8dwiV31TN+yIk+Mdm2Eh1vUsOqKZ3b66pWeEzARjQcYIh0O2KiNr0vKhzI
OWNgEH0/HCV55E3QRZ3YB+4K86JawLGQO1d0BwtpdSVTOzfVMHeNkmkY6wfQI/XDtMCcE7E9/GsZ
wrKMPrGe9av9dvaqaZi4HBuQuyZcPPJXk0EpyZGzeovOlg+I53l4keQpFRXKboD2I74/a7IKSBGL
nWNocy9ucLUnulCsPtP9y2HN2vm/HLeJm0/mlnb3zXEmYiNR4wm9EdWAEIq/0TlN3rIkomr2sTKW
kXu5wm3wwjsj7W3xKmnCA1GccxkfSaLCIfoG1ZYse8W98N33jsxJVB5jHp2xCnJGrH7WtKeBnrFR
hr4jTwQPfKqj373fbtsp3ox3cQ/0vnjS69cSgp1Mjr1cJN4YgeViA3Rd69xsymWiHAowSgLj9JIH
qARKLj2wy4JKNGwIFL1vfi8RPSJtH8gKL99gqPeIT44dzK1usHAMt8yUc4Ro+GNWcFRDBKNzL66+
rPy8+gy/VcNeMMG2iAiNRYILQdLMmOKsR+Tle7mTHI67PgPPG3SnDOXP5z4PBrafiPOiDoKXkPHa
6D3evpsS/X91Jhn877vUiphOWT7rrPMNxQGUaXB94mkBApcfjj/CRyJjfO4BocDaoRIxcj95wqJN
8UtvbEaYfNYvTwGMZrNAWZnZW0RJSAFzcfSSskMbzVKepSIWzSTg8v5mCl978PPZjXdks5MG01rj
VVNshAoGEPqK1OHh/c5VZFH9G+frZjIluEcHYCHbeGaQld95l4ZYVSzjkTDWJQ2SM+7Czyf1hs6P
u6ilMkulIArL5rfbOO6Z/SraDOuGFXPIWMEE7jn3nnGfF/axd6QL+Pk8oFNVEYf5gAI8bywufWW+
fM0ahy0PFW/I7mOiAcx7Q5/ttc2d+wyXTEky1Tp2Hqqi9PtauGXFcxXD87/3Wy97yYNyYgFkN0gC
Ar1IPkbnvx/GJwJKiG5740saqBDuRStpYVMRr5D1kCKvnNn0DyDVM9jAsXk9JdzxvsoRvS6ZFzUe
LurTqoJDucNLFpOXEItvlYBVcdXla766Z0iOV86QTZCQ2WaVn64D6vxhdxNnfnpvaO9gKCOVo533
HMQ2bCmaX2tD6o5+a7ElFkA5RZkSeU/66Er+GTq5i/LevevpPMYMMxgmgVT77YKSSPK1cO6UHYHG
ZoUOn3S7EgHrJL5prRleeAQ49C/bEmMBE9OS7oH6PmABwcnm52kK1Es6ltBIjyrvQ1J3vaKV3leY
9qRx+WM=
`pragma protect end_protected
