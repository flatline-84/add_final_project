-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
umFNCULdhUfXIayUhly9H5Yfqt7cIriA1XeVns77V/Nt80HqUAXICJqbUsCY6tuj31gw5AUjddWa
a6frnFSezOYKKpDomCYYPohf1EKeLJnqQ3+KA1OXiOIINzyXnLe5xgMeMITCoyE9ftu7TDb5aV32
SEXivU8eu3mTFNiwIdeYGQv/RDGcYUAgO0iTE78LU9nJUZa5d1manUhUZRoz+XoCYrFzW3Js54i1
VjiZNi5D8hqBKJo8S261Z6uYzxvRRkfd5rf8O34eIgq2gL9MIvhacSKn/4jGtrjqRAoyLGLxLaBI
ELL4MC7hcduR7ZtXxfROlDOQy5xU9I3kbLZuEw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25280)
`protect data_block
kvgj+kHIsBiczRftqgTzRmQbxgsAkAfvHI+PpAg9CvGHIVkeb6J75Govil7s3NJC9lCKNaPXQImT
23EFAd4NW6egPSxwgsTtV19r15/qudSTGWlcdTKg3cjQ4gv8qcgR69h9/cH4EFcQ0syIzhIDiW/4
Rkm4c7n/IteAU1pduwcba3jOcfirLAWRipPYMa3LpFPQCQQfSMnRGbygpNmQdkaXMu55EauYiU1M
wFYYB43aX4AhXK915qZ2PArdjueiaiom5RvAxE/OaPCUbiWugLChZanBwE7s1d3JgmuOwgr4R4O7
RRrLAykGMYr27Oepj/jOEAe72e869524HKn93886mb9+yk23ducLuIRp30z/80pmLQlKqKdO6F6c
eEXm3gz1dTHVorfOClPwfqmb8QiTcRBTZAPvjJPFcSM4yC+vD9Be0OozWTMc8FVlvtkeh4opjbKN
FmagB+B80aOn1hbW4Pck4qYcH+g5D6v0M+nmnzZ0llFL72IHVT3iiwad5keyECM3p5HNdYDN5vZc
+lAm6u5pUdagAjJjAgqMqBQ8o9vI8qXFZdqT5gE3t+tSXOrpUbOU8FKtuCehMuWP5ZWaGPOHgrkm
qvhW0xf45agOqiF1xQUS0M5d/1BoRWhWy9BZlPDM/a60s2TSmNYIVZM7WEfODVM1Ya/ISrmIvqlV
m/lIf/UJSUw0QCREMaME+96X4rQ7/NOVh3A9QNIKdwC9FVzBfsqJA+k7CHZ4JVPqPJpWgsa+XzP+
0BOMoeincNHMMRcjMfWFObyX6OHMKt3arrrEa6QyYK3maQi48GuMaRlk8+IhKW1DGiZlR7JZxvN7
LxFkAG9gTMKuXgKOFVGDelraT8tulFJmoE6EJ/TQyHuGIUZSkWhZNzaXaqj1hXd8azzd6Ujxk8ox
0rVcz5IEeTZNJ4nmKSMMQnVyxD5BY0m2LUG5Z3LrBVO6lvLnKsL9QLK7ly07fQICsm+2fzdKoa4/
mbNToRXWwFQr7SchAzEl0BBk6cYqTz2nN43eQqvh7uHcknXNBVKdwT5aGUPpHnYemSKsZTjUa1D0
A006FR7CIPqxC7f9+t5fOmSVmhvoDm5la9NyApCEy3nCU6szssG7m+zRU25D8p03/yP0VKuZHQJS
+gioHf9wXvguY2kul/nePwoXzJinV9CKqohrUpAYx1KTSQbIaWdP8gLNf+IHyPYI/DlWcmzrn9ZW
Bz98yac1ADWjKoLdt1Mighm4BIhRZAH6WJKFfARVo2O0U2qF7lWm1MPhheysgBeHLDUl1E/L4SWA
1o0OXIO8CvYkN8uYw21FwayxxDsAbT0ftDb0OdFkQTSm9tf/VQNKewzZ16aijf0OltyPRolgl3ap
yEBnr05BWJ/8CyUI1qOATxdR2DJFOM/I3t5cCg3/XR00RCQEz9yvM1Cw02H9aKsTSkrjGn1oYrzz
vXh8rMITzL9h1s0i0fLOHPBjj6zq9N0UoZeMjk6VRVfUib5mYVlP6boYCm0/HzoYgej0V1jMuhEm
CvKJQmvoW9u5q8Gj/suD832tqobriHAs6jGNluTxA/Q4Xp2o2V9U9zl3jUKvnRcakH43XZeMEAGL
Uy5oBpB7hPnqjr23Z6UQKMaTs99LU/nHsFmK3ESLBb4gew9xm6lpeqCR5kqw9dH0lqbroHq+zRKJ
3LdSGK2q/Bsn+5YqXLkyVNpSRzUWrX9ZggnMjFgkRIjTH2jt4tMRoYmTUKyN4bea6M3v7h5fFCkL
oja9Z1x1nz5ZS/7qFKFGZsXKvxzVn/6kALuFHj7nGxK7LEKuilo//ZNuQe1FDYthBhxrO4W9bkeJ
Ey68RmAQrZYBUpE0WHVL5K9iSYq8H0K8Tc8+Anizqu2IkRnsZESCYH9khxK/plZ4t3YbW0s9mCzt
mYd1R3eK6lkPWJJtGe1EhMUKHQaf/lyKQdSYDpaQFGuFkbN12zkfLSegi6ecnLAlLLzakrNzGEsj
+ToWTbLTpG6ImVkS2zYtjRPPXRnfuwQQLiHsitq9ZS65olUfVmdN40cF28dnMgsUN22yBKB0iswL
DtkZ5hhLtw6rtlejRerLTYwT9Ae2you0lpja8gv3gfqpmFH/9wZGc2etMqtcJofJT64x1Rh9BIoi
AFSaPASq7xh8Nc7eNxzXHYGYkNwotGBuJ8bTz/sIAwsYyfIKi2LrYydFuro+GRoc1/hhDOb7DeEC
S+kjZmJlWqV43TxtNjxiBQPWkX1NSLw+GWNaakaQhXvDNOTIrrLtAexZ/m0SNFrQ8jET57iymxnb
vlHeDKY8zwHJXn78fzczYZr6DXCJEQ7h6oIFx9FZ4J4twH6VjAnaFz8PavrIsB21CN6QvtLC9ZNx
IcujqJDa6GGOGUbQFxJUdz9Xsf7frcaRVjpLtkiLomu86FZNb4c9m/f1wH986c3GwD2DpObQjq+G
FaxE292bkNtEyIx1BN19QLE1ckY8WHXSo3rlpjhXDA7aItT4hITBese9+L09UYIwb2T19L9JhvJr
np7UBf5oiARcu6kXFWC1jvIdgvXqRLVumWb0TrH5mwR1wpFLzfRAhoM1NqXiWUZgNcRWI5UJYXFS
23gCjnCyjBvVZ3EffvU5tMpKzyJJFN0VmdAQF4CeR/XZGTg+uBDPDfBRRzeFMd+TgGKbV/zLA7oR
SUwCiGvruBxK/ZolPYklLoJ5pEH8zZ+I3HtoTFxqdApeVsKPzktYjYqht9ih4z1JVBn4sjNeLWGr
9wPKXlQdE1p9Tm4AtJbTNDodTq33S+HUdWaTS9CdtXyJ0VzR25dAXRSyjYYblTm5T6/CeEIRiqPv
xoBglZBsrhYi4Vr6OBOpG8BMAzHX8SzKAmH8aqwJAFdgKCGNqKnENOYyRse4OTeXtBvnT9uBoN/z
e8VVQz70KI9NlQorYbQA/qDdc/3Ff/0/fM34/WALJVZnI77UhYd1qxKxhqHE1ZIU/yTO7GEwQxtw
cfsib8LbIE+zyJgXhi0wOFE/Esy4O6X6KnaACOReVJJfAOpnZV08Mb49XsxlDJBVCrQtiTdMHZ0c
CCT69wzGlW8xATUY113uxN5AYxZshes378thySsvVC4IRi8ajzg24iq37HFah8eAJn5JD6hjq69Z
cZ4RGSHfAmL6B54h110m8vHhGZVvmzn8D6bqPhqNaT/RvjbGXIS/gV+BsX0A7z7SDuHLkk4O0eRQ
JxulrROOpbV5cMB9z2RPt7enfHTgmPS2NBP5/+eCG8RpXXZuZtfqryjLGIGmfSK4uk6RTFGof3rH
DaeOT3tq/rie/+bTByoJ0eSuBUFY7tXjFdyv2bh1cbqFtwOnTcuRyBlNV9XgTyHoRiFjBwLq6mvW
f3DjVROB43FRr3oo4aPfKg07Uj1AbwRtlVF+az4WP+GXtQuU6BhVfkfhQ1zXOGzAhJiC8qhAVeyz
I/uqICkN2xSYkJIC7cum/eSzSd+/MbxG7mMrf8cT2lGXcnUGkt/W0zYljM/Xme20xlvVg1lFawvH
VXxVbQNWlWnHC9N/BG2n7Gw7KE8mMcfIQ8IvEwXA8OjFYs6k3cm+EbBowkZnqXzpiL5xPfiT+8ty
j8iCDIl7kLm4FXMlfmCGQz9vlk9wszBxP5wBoblaxla8nTk9iX3kw1V4UwnPS+9oHqnammdlR7dX
kyw/BzG7yFKnfYGe293jH5/plwoNekrysTKunxUw+3CTwj5O1i0XtEgJ5ewNwYAGXau2qToE+6nQ
6avdPRtZCRGY/YTuzOWwRin/52595lxi0CY3FVw9S8PLslHRQ8gNxiyVn9BGxgSN6dIOIV74h/3X
6MPWF/M+2eaYplxWzHOFyDFPgH6V3dTiM3bD+XZjlq5xlcOTrDtZW1VnBmYuO23SiZhDhioi5mph
4IszkniuQPEMKkGKoLk6f3JuueuMrt+P2uQafYpNz1tpU2XXnHQyT7PhgcMx416czgPZ3M731yg0
7xCtEKpCVGdYvd3xbuaBszoA95t8Df5XmHh1FUG6ZggoJ2Zy/uP/B3wkqBPoOyxihh3sNRQ8zYbt
Y8vThAhldY7egL0h0bJoZ3rHmRu9UJzSxZdTKwdrveBJhiyNABaXC8HoQMoJBDEQ4fSULmyw5bQI
MccKZBY1tDly+n7EFDZnJToeJdU7sp3lbOVBZynO7J6hCoNdA08upy0rQ6asHGEV8Ou6rSgKS/+p
iryc/Km9DUiu4PitkPAE5xV71DwKuA8/Ze5vS+BfeKFwgHKsuKEQ1TJQW8RuAUt0Y4CvuzVfA1qN
yUQXynO60ClRbbCmDNdYRcCPylH4bKJ8ip02PCbU+aVEk71JspiRzqDcKbUdQolt3r06bPK7iBcy
JtAN8adM90w3BBTtDRrLY5JcW5Ios5/kZmQx04kGHkcfH3pZoPb1vqdCXO7/I+nONiFEm7hOR4jm
exHXEk+ohPHhos2blPusuxDjEvfTy/V0it+OEvxcWRtQQwAiKgERcR0Jh8zT9PkAEpHb36jTMLpp
dSy9RDgMopaEfecA/YTdPUMbcwAQumCHZ9834GCgangktN/jHvxU1mdKKrRii5ktLiMmW2+v7/50
dA1dhsU//cRNmSoj1yqG7uo/HnEooCiyHsKgYvleDUC1uQJC3QRiDPhWDuAIdAesrHi5GL1yXfpi
1FV5RbCxvqkDp9WS1KP8AliuoCI0nakuwJ7kUguL9rGBsEOrsxGOllS8pTALHFDrB4K+EPo3nM9O
1IFFKRq6IMJWYLpaSwMUdLu5epqQwipIrrU4DSkdICmVllLToc1fziQNXiYTtYxtlzb/Jfceqsmu
z+tF6lR5oArC3MnBDojm+cDyO90xsdauHaZvLvp3S991nozlwgx+ZW6qc6s8XaOspPUVUPq159hs
e5wlRZRMu4jtPszYidTK6y7dGwlAyWzb29TRd3jf6ma7KKOIDMRdRTy87nw/ck+528MBOmilunXO
rM3ZHq8DTUh6g6CXqt2L5uWsdBDLem+YgHCUj1UFK/AungoyVowo100HQY86n2nBOCdKBbWgTIxi
vUJG/HhJ+PIjP9FH1yEg9jbOuPpcao5oODK5FYMjhZGJug+WaIsWe4HoxlvUUb13BdvPY5IEheIB
+O6VCIETzVLSJXz0g0fAsubKiRCpgQNAfnrbJNnKN7jJDz5SZkk6gFwEfZas2fVnadB3fYpXYEA7
FZo0c62kexiWwI8Uzxhw8Gev4f5j74Bcl7/vBjQlVfj8OwoZc1LZoblZNxqMdvYi8Dy9KIMHXv6/
XBhC1Pp6/zq4ltY+gJK1w66UVCEtioCz65zNp0st5gVXIM0FxMD6TqN+9QnIVul2vaMaWYPfmDJa
q5X0TBGBJ3gwlKnvSBpTkgz/P8MreqwGWBVcF/ARWrAaU4RXfiaXPgAiraTFt+KMPsKTeakK6pas
rCIb8aKMya4EjQBf+jcWAYguTPCH0auQuJFM1wwc8Q43VOEVBzkVTDSXQ4VH7HNcj7ntpBS8A+8s
tT2SieMIyoz6SSIeFZl0xgn0Ad+3EW5M+tz+MdFqAkNIC0NcrKgJTgxYjCAwcUIg0ul4ISIYvr6q
1PFPc2Fdw8MYf07yVUtlA7RA+XZefFq9o8ME+W80aIcFXVCPEZqIm0Ip0uv0BrEFq+KIgYzeWPSa
ZNdSKErJAhpTtSeP/7EySoFKHkxCX0vKym10v+1odrlf6sfGr2+kw3Ud1ADWLnFgl/0kisaQ4gCR
oK/UsM6/zE8puuBAWOFFSXNx6ifNrMznXO5Og2HMrzCz4B1KduqCTLhe1UsIxcIUsIVTriE9ITlU
dAN0YS6NsnSmlc3DmMu5qV6jU4ffFbtQzxi1ks5G2/EQiKpRWpvwC9zryEiV5oXYXV/t4a5iv6To
HloIn2NM2oYDyG2s1qIQXEm169Fm5GJBrr8Ck4eKrEcLwLCdqtcwIWthZLTRpkdrNVPr8VONHZ+Z
1lWEKedjBYzeO8WH3qCzQyWB69BXFvOZidxDs6TW2jHSbWrUvhglVRU2gKFWu8keo0dHjLkruEin
aa1YtitqSInxAhPfQKdILIVHDo9bvVu8AaAf+WW412M0x5DL7sHEe9qkiFnQg3u6eOKyC5cFv9w/
vAr0DQF0FH+jyhXe6IWbptWNjQ4AL6jpKweOI6TxG6a0oRvHHzaw+5KOKkmWzRehoLDK+JIHfq0F
pwJp2g/xjHBe6bTAiV9mQ8r5xYTi5SeN6fnU13jaFQAGO3dD9Y8wMHdA27iGV6LCx36IW2MXMTzH
En69uciB+vPXJv+MCIrvILvy45d4U2L0h1nXEalkKWaAymN45Zcay4fmm/V2aIrRLZDKiS5ub7jk
KJ4/eEQrDs/JRiNgIza0H9bLRdILIAbIscKEL/DEG9XO/gC8LF2hqsUifP2DLc95gNhpXiTJYYaZ
edn8QPSr+KidoRTCHwNAZHWVP4uDqEmMjON/rhmxaHcTrwFuiKIi0Rluyr9TdrnH3ApAYV8sZ96K
/IuWsdLT1Sx8VHWe79da1CByA/QvrHQaOnbNOVdwPF3LL8nvRSqPLTQ5jSWJuuD0HvCwNSpXq8Js
4i29o6NF2S6Db9gc1XCFjF7ZL/ZoA0G7uiCkUb86pdcffg9Bcf1GjLkiaRJIHGdilfbnzZYZwCH8
0o0yFoit+DwGCiaVFnuYIwAWSovFagwx2HTIZ+qJUA+8NB+h2eUBel2ha0JZDkV8msMvHDtiAP5O
AcOIISyfFHmNj/otQtoVOaES17VwnjgK/ulo+NYDRL4RMsdgYnCJ+Z+xN6ZM3MtF9dt1/tBL1zxs
oX/59hBKSDVAsXPpW7QmDk8G2pwJyoRVaKqnmAEmAjwbrFRwRV4NkbKcNyn0RXo784gp4gssFZM5
l49gS/cRcZxkCR7TMysjV/LTOkm/Wdbw0KSSYbiCzGLtWiFCxwThlqPIL5j+GYrzV2UmaGR4/ylX
TfSD/EWn6mOV2j0z8+79Y5Uy8A6FIc9g7xfQ8Pp3aQT9d2VPsmShMogtNj5Ufdd/4/EuxHuGUInX
v23EiA5VEcGdZsuxDRHepZlKNl2GGV0kCsvf///tV3CRBOcLCVGQiDAKZ4T5x60UIZOoCwGfY5wz
7tI5Iu6XTYsmdfG+/EQnUe+jHitniIFt4r7X+9tN5vE+Z12RZl2JJbY3L0Q/7ef+WreORXVzpIVk
SgujfjBIFA7uhK03pCXqpxU05UFKHWu0qW+axKwHQ9fXmQ+6Ahy/00ytKdHesaKgXRQk+duL4SRo
LtKsPVP05OV+Tu0/T7gNU80SIeLl+h4002Y/wzswyo3+kQo7L3v69/dNUJ7QE/RBR3hqkwmeBlEp
g42a/4dmvRqGoqbzRAyar2itgaSaVK5ebR4IFIb4324Rhxb96lY0Je1oOHmi0rIAWrkuBnNg5N+2
PUVt9WTqBi9Zcdtv5cXJ+vNvtaGnuo7G/BYxIbjFRv9Ni0OQlyi3fMfu3ZTPzgN3pT+fCwDWazRN
lFYxPFhlkm4pFeukwtPEg9Db2wsFnrjOYsgqrqJ8HsyB288hak33Qpuu23fhI6J5ubfqvBAAl3j9
7t7ta3zoBVIsVh96lAUMfaJXhEWaBW5L1qlJ3kPUVB0Xw4lYlX8HAq2F719cl58znuwiuyjM5a83
U5cAbYZanMVnJkjeI3u6V64fSuDcJigU3e494o6LKQWyPhcja/XOmY+IbyVhzl/jw7NIs+/fni0L
gowI+X8nOTEVYRFocCF/kQUP8cbqsqWCQGtG3yluU9G+8LKIKmO3+owDrwdTPagc26Y7VZTyx2gv
/oLV7r555O6vRF3MF4LijlNL56XESqki5LU6U3K8jXxqgdWFmt6qHi3atiwuIYh2WXcnUYvY2TN5
wkqKV8qA7fGwReXu07ZAOpJzhpDXc21pY4Xj4kAas07rBep5VXYTW90WBYdR4XQho7XsoveO5xTA
B7Vjy9jsMusefaH2yOmklNU8lu/oc2WNuS2lOu3cJVWJ1hlq2qnKLXEXSzA0dCtY7+tVEwthqsiF
pTPuxX7ip0MU8aI9Cx5nlKv2u6m1bqFgLYx/NN8Gcdi2FSNZ0kUoGsB9W8URN3gnSj4Uy7xoB6jA
M+RvrVoSzZCDoN8JgS90bQwjWNY1S7p8jvSnIoXy7+yQgQeAL4NMfsuVQ5jzfT+kpuQzCoQYg7rq
i73VP6NZoUhmxKs4QkoFK5tsHb2Yh6+k0WAkSrtkK6kiYpuWGB5HTYr1bvOviPSAZGNX2MOFV8Ss
NCdJx7e9dSYTVxP4yo7OwS/kO+JLvtZ+Nf1/FgEanBAiVkm05Ni/Wbv4qcadRis0FBXRUqgmhwyH
4tVJL5iImkAdIwiauXBMbTxchcKi0Q/85/hMIWfV9LjXTrumryRs0E0F+L4rHBn0EkEjXyVTzwg4
Yui5pfqsnZLcrqf2uf8kAZ/ysuY/Dr/uzUh3mbz2JcK+DB8rI9cT3sj276wOv14hkRb4alPF4G7Z
b3uXUILKlVJh21hhOigtufjXtC4LkXL5RMkybydzT91kLK6LkkR6396iWrJOtHBhMIOykWgvUvFM
Wk00lgmPC9vstseMqOogh6mMyj2GrlM6Z536ehnHV6fkCImwfSYqdxr19v+r/uNZId1Qb6pGbMdf
pB4X+dQTEtgCKKX0uEtTdtC1Mnd6CbjNXIKMs2kMV8+6kFse5tJkyMDV4vs+rSpIJWOCK1Eu4Jrq
4DGOwLnrDYRzw/a/uQySGgrGwpMkP9h8eWbrT45WcPe+PDOL1sOfAb/svaLqRaWxeyAUOryVxkqF
MVhBmuz7Icio77AL4pnvyeVNibFkAfpuU+AKK9iwLeh5UzplXCTeCV7aPZHHZEQav6JRr1lhw77p
E+v8bl0+L9k4vnUZwGPhkgY42dWWj5ZfRBcCCjT0pY53ZMBJMzhEKk6cu2L6DKFi3gotOJfYADTl
TX7E1Ot4rz4CrCh5gyd9VaMsTpZZOsjkwosuygt217tNTFHsOli0alQue1/IlPeKEWZZZrGCxRkY
Jt3Iiz2w7nvl1qcvRLvdPV8Ga2O3ov8Ix4K4zASwEd1u/nRthm16Sg3+1JuaCgnpDH/ZDON2d5PZ
6E0zXk5gudT2QuIn6Uf3FWJZ1QPrlH65qeMfxSNMpR+A42yQCM/ex5iMVXHbHC4BaoIyrsKzafs1
js71gsYPj6AJYyX0Lt+czk0TKIsuP6bEaLQRtH17rJ1qnb0h6YlX7qpJjlNI3XnPV48v6InX+q0+
KCu7OEbV8DzT3RZwbQ1vKDyUD1qkCAf/QzjG3KNKdzjg7KN57k0JAVptvRq/bBrS9K6Cve3S+H9d
bQ+Z0pj0H/+Ze5JdbsSFVpWGgnZSfVWq7VjGEr4uYZrK9LjcJyDdo2Iv54I6UfAncf3pTuAKv+E5
QsuGJtiTCTzuNEqY4fN/KMEy+WTsL7DJ5InHi4EgDgw1yfYe8WHq1fPxL3KYYo3RzXSgl4FnbIJ+
mhBO3eitGMillO3kKTcQ1eZq/P4OiA2ywq9AxmEYJ7PdpNvtxoQ+g47sCNbSezosMKOuLHmcRZbZ
en1LhPlm3woWV0Yy77qa+li9s4tirQNSJ08fgO5+m9Z8gK+uBVj8cjT8a4dYv28oL/LCFVMEKOTm
fC+c/7Qd7JV7fj0mur/bZ1Fcr+YqL5bhjTNjKwe5m68RogpXtJKTu/y/pRXxaQa1Q+UrhbDMIHnZ
HB9u4uXfLUW7PMK4OHaazNWNhfqjTbiFkiPfBlNf4V7UKzKnlaV2VyQvJKEEj7l/itQmNbDAo9qe
tca3jsO6Zyj4J5pBtiJMOna6XOFlIeVa+uFDR6RykiGPW5fXne54KX/CxW3Mi1d7IH7pfqvo781j
CpuNflqq6aOXzBc2JT2QVVtmmAJKB2fUT4FYgdevGYnRnvuSRmBSKkKcfHnsv+TERDVT01UoHInB
f0R6ojGbj6FwLSTcUtm4lDaQ60Yn4GjMwhjCqr5T+Y0Zvl3ZzHgVo8UHZlZTOeUGMelnkkF5mLmb
yK9EjVHIrVjeaHx2VhcWnexDultNK6a8QvAoNfkoECpXhs8EzIkBUXOcnynCAN4MvAUpn7m00wLV
9DPNZZejRJq5S5M//bf9M93NHUeHKTnZCTY6JgRsiyCtxE2WWu+e0VDz1HG+/tNuMarUSP2wtgM9
0Q7KfwLaws8RzaBasrdxFFkaEIo62b9cdaE5FQ5PDEujwdSWkQayFTbkZj+ocWm9KPnBXz2YidFb
k7jKKbl7oPaM5yWloHUDQ4HHVDK4KsNVm69PjRmpcBNDLmxUEpn+mRg1SF6JnfY3HLd5vlQJq5eR
O5ALBDTofAQ6Pc/crIKG2sJurfwSpXwvt9V7rdONUAo7Kp8uOhIuL/SSX12bN2ax0OgpYbVacyrf
f5+/oxZPHOm5jrSSPITQNeBRAokLMesYMmEapZJEB1CeV1X0d/1v8LZFFJDjJll89MnGGtEcv40b
WN+Ox4CIzOgAfKV7t3gEpPQ7bE4id1Fa4TXgffLkUWoM4BJbEjfzjXyZTLAuqIOpOgYHdJDL3tpq
ivpU290rEOiNoM0Eq1fYpcsP7JtvOFH7d7Emoj1KkfLuikZxo9V/wqpPbtTvgz+fqTRvlXq3a5IZ
XKj1miZhQq+ZQK2EBsPyUyZG47kNCTiOUW0suBv7MWh+8P6WD3nZl2CwGdTAhehqbPrbm8Fi6InK
IhkcEWZGs2bvA5b/CYO7XgufnsqUIRl0DFFV1j4Q48J4wgCoywKBxCQp5rge00UzC5GMnDw+Vmk+
RMYO7T6RyO9zyQdHV/b9wyDelJWyhgMyP1j2Ms1TItD3I21aBMJGeiKpKT13N+nr670mL/t5FgGb
diVXw5EbmN378dChot8ZDLNLILL9xFk9FnwkrSjgN852pJlQyY8CIu6x7GY6z+6E93yPMFeG6hnW
AFbnSMRtSH9y+aZXeIK6uIYw0rH2i7qglBWU/DJskjw6KcUvpJzcOymeNOPPqRgOl9Cgg2NAaKWL
Ymgn31w9ugyf1gO2XB4M7w2z4baYepD5J+9WLN7t9DtaKx6wJ1g1tLcDwmPF1gUXw7gfVgLH/xMk
LQH1zmdeTKyJkN8KKt9EpaWOBgluwTpYgWavz9fAHtdNGvLPlfjlS9dTRh7+5nkpnkaW3kcSA8S9
v5btUONS1Fl29/ZWDxpGZJ8iwt3qInMO0jk/mxX8rlVFt05vMxkx+2f/Ns0NI4ivocVwVJ+ep5nl
zw/gL1t0LgwyhJ4x9hWYF6dqNxvgq6cqBbOslnzsWChTi+PvObN5vUOsBPdlRi7bb8X0va+1u25h
96kvLaMe/VizOJXhRZc46EErS42dyu3mMjPOXlc64R5vyZu5StvcrbzRzGr9wPiif0clV+SSZlNH
nOm75mAXlD77p0wXG9b+FL4CBXg2HRunZhd7WB8Pg4qTd92dqlJXZ1rc7kg/2ABSVeTapQNwy3Gg
zLtkPZU5bHiA3L5dfTQsb80Mzw9MODvqtfz3nhC/FJUx+l0RAR2T4u6PNI9IWGSp3x2+wIboiOGD
oBDMo53aKzfsH5hHvhZS9FX68q8KO9yadsMx92SSh6KiJ7SNAMKpZYM99kt3qAkCFyznaCAdUaGC
f6nngMv3PfigsslyyR9h7i6u/vwlnBwa+ddVOsjdfRglD2QGrQ5Nah8ZEA3v5ZSLc+S/A5rSSCsJ
kMXidD3FQe9ysAu//zASDKwgWZKl5DcvHMFey9glGdXrLq3Rxt4ArIL31cqGl73EtFrqPfVO4xZN
ydUX+CngpN6tVSypEMYR6L3TSN9yNSes1bMtX8ji1Ku0UKz4Ts4OSwrIl6nfE1ExUrnnCroxvOuT
Ht0SL4IgBkldlZqgOdBY03MtJJqlwdkEkKcNkRlmMBgWuOR5Hp/bBQPpGxG+qalm+mVlzl8DqXyg
4kYS8Sy0pylsVFAek9adSwFxdKbWP4n9Ne/lCdKmYE7eYixak6LTh2Leeg7Py9VQYMTtiAy66usB
hisV6JlhOPcIOQLfkugxJG3x2Fzt8l1KFwkf6p2hByupCAsOy0sWl0u+CnjyZAbpowkgh4Vjgzpc
Bw3XGhVosXA6t0zxX046G5mOQ6YnPpKT6lIeVBMRyVK9KDepMo0z0yujV336Lhd36ILSYkwFBm4b
bcR6NlIa6xan0n0ZQjM0jhH7A/qWUG0VhZiyoLCBPKn9espEQGAiKdlDWXsrBmjTn/5y9H9hwCFZ
7rZwSOq8vmrYhDGYddcxfODc3rseel2iAK9DLai2G+pL22x3OxYjTLpFE99noPECF4t0UXKV+A24
F+gbcKUf8rAYhwUa4MAWjf/gFNX9J4oh8TzIn+8yPVNfrgHPs0+eP56CeYBAmj78N1+zStMvAuEn
A0wn4wWlT+zMyjMQ/qGiTJmIiFJgGpnuFOISyg2o28Vswq65LwP/NWGGYOtDU4IH69+eziDSG38c
O9zFEyvPDnH7lWIe9PKx6VCliekRDniTIa6of+l24wPrKKLgMVeG3pKKsOfHbgGf0inGGaPCpWLq
VEYFP7nEAqW1ToLbnVlqXJ0ARLMh9ux9kisdOQREahVKYcURcXkK8KE3eDZhXaWQM2u83N8YbeKj
XK6QaKedXQRnxCVgBNbgXq7fnOg80Zic6ZWlfIRF9lMH7UMLLCczCiBmkLzy1Xz3eOBLhrlC/F7y
HSzRC7McigRJeJmhqN8fZiVoKfX+izscvQXCa4WWBoUcJ1GjRuSU8ATpfbZiw3Ma339H4v8Hu3eS
wrEw7DT6t0mqzQTZUYE9+2XA3oxrs3XH8PBKLxDZD3eN1WBQbzpc1dtXgqsAJNlxMGbiwvCldxDY
9xG/nN3io3sf5hoz1ItFWyi0EfgqxFarNtVAjkUwroiLlJxnIszQx5Jfaz9hQ3O8nOKraJnHnlya
eQSaH5PefTAaONT998JzbfUTraCY4KR7iu6GExIxYkC+DconBSd5oKQ8gxXW1SAR04xRi2z98yDb
KHeIC9yc7LEc/YuKdYmZNzgxxDumk2ZbJvZ6q1beOPmnCCNpDzlkgOKgJikRhNPWyj39j9tfhvit
MFXExrsQc8kQYRybHAR6MTkigrt2urW5rdNSPeoAC7BBfUG99VDyD+69pVNDAYqbGsHmDD+BmST9
C5wsgx9iwgR8nc8kKHIoXMnIrMir1nFPtTDBQHtQpTZ6FK833s5puwXHqClcnpKeIGrDsIq3uDki
svNq6woz8DWPwPDdLWp1xK4Uf2mr8IOxC40ESZHPrHbDnt445HmIFIHPTmjjaZOV8E5FPxtVc49K
BX9ttXueBqAbvjDC1/9Lvi5EPrYxJjWI50HA/U4IEGl4RxS2BilVQLUqnIMtWFp0LU9obZOeG8wd
LGarKEI3i93ThrWhav1Ok0kn0sMIzVAsF5tru05CQ9V5Mqp4P1OKkuWpbVLx/xCku/aWzsjRdNNN
/PS8oIBkbGUblUp5RW2VxMwqcERj14c7sa3KYuaX5U3rHFjIZrhYFItGvY0sz1EgRvPZ2Ch6VwD3
1uM9EJVsa4gJbeF+04Uho8zPX+qcQD0B39UaiQCPQrInsGuKwuFIDg6+2GXe3shT327fGPb2HvuO
VhyijhFa45FYiFA7oFXBaxqHEyuTyBPmKKCyW5k52E4XQn1Vo0dHws+etwZHqa5pKK1YgkS/BphS
FGRBELQ+Ud4GTq1Y2ounTf5l62e1h1wrAZ9aYRppjodxdiueVIP2Y6NAgj9JRomRA29qbOomtJke
k7Mqh8Itx5dnqn2//xF7SN8khTXAUQlJVpycdMJAIyhOaVjYYh0fySiQS8nclZSyKIKqncI7d9VL
cc9zrgnI6unnxiM2LHNF0gZDlRf6plToHoD7i8elq74M7wevggAxxTgbs3moPRZpttlIUZrT0MFY
7xJ0qfFT8AY1bGsMMLEYjpUmRyMMCeBA2ZMFMKpquwJ+TZlvgs/a0MgaFp+N1IYLjt1I403ZkdcQ
zNShOF6nfzVzwza03FSUzfjMoIDkHhcnLyAUCXQLNkP7Xdpf6/uQY24A74rX8jrO18lFgS/xt/IJ
lauWrUNNRI+hVOjOcx+28Elko4EDa7EyyXHgxU6YAwmC22nZtiqcVhbecaCJDmDB2cfdU6H1xU6z
fMzGKp+N5HrQBG8s0SScNrhuojkSdwMo3jX3w/0veULo1QqCxNbvab1blh0nR0/VFhP3U9lFYpdT
OMyuFWA4N3gcbtdtGd19iJUFDAqCdBgfxI9HBgQ6eB1NWRHg3F5wD+fFXNeKgCTFOUvXyFitCUGp
C83nKPh+edK1MoDBUwsdqpPDi32qGmZdBfyUlW7ZpcmA54klkhHUJSMcwlTw5vdlMjeEqbeYiaia
/KVoxWJzw3K+Ff+dstRZjOlaZiiKK1gWPqaAV0/VwojBHgh1/ChMx8tUNryhgBjFBiPis/JxzVuL
8s6sKK3IA+oWMY2HD8VVq61If52TvJMAlKZHI8ZcpLo0V+J0n7rzQRA2TIbZns2p+HoHm0sUqJMG
ZujJEel38nTNYelqJlTonnOQCh/n3scgbR1+1qDhuONf7MiC5Q3ChyviIeffiC6PMmAc3/p4THxj
qtoLroCmWYahocVnSFarDQxzD1XKrW0DWgeE8tD3Mb0rKWKe7zAdghzlvRqMDqvSI+g2sB2va7C0
jrWWBqq/gfMkYzsz+XV3u2l04NnbkBeKFhjrjjK2/Noz+mCRtOSuzFFyTSZAUkwe3MgEvOYiryUJ
X7kDFT+QazudzGu9aBZKyd9Q7YzcyiY24gXOTj6324wql/ZJ7B7vkFeQIHBEmtCuyq8gRkqHDaE9
epUp7whNOT1+CQnq4ZeAm6u2Ysb8occJyIzNiclM1NM5/CI++ORdiPhlGUM5+bYRyeiaM9S9jjpg
ww2ZL48/e4IpPpdOv3pPBxkzfTbCldi4c8YK5O2jifTPQF4BzaCD+M+mf5lYrU3skChqYYWhCqAr
DYtB9tJ5q7bz9YbEgpbFH4g7TatjdpZoj8YXDO8JTE+oqr3XGRbua/aGY3eo//VDQCTeiv/97zE/
ZUYYFz7+kBjokP57CgY0rBviNU/Mp/myiGeHljmHqscfKUHC7ue4vj+rUgHEZPsMEATMN1SxK3aR
OVP8mDmPe/63+kNk5+AT0nKSmD7csLPhxIpJU2LstqYJpU+qDQyeBVVoYg5wl2kQIkfD+W3wMjxj
k0AzSaQrbRHFWTSQfttYiYWPuvUjWMfdm31Qh+dOl+FlGeg5IlWeSh4S5qEmWu1HCDGzjq9sl+oR
vX9H/dDoR/WrEEBbCR8EYFdobxW7b/pJ7IgP8xHR6s3jFnKNNgLD5pytZ56hIdKDPORbhHoVlPD/
99Hlm5Z+kWnDwwGV4Q6rLPf6ys9AVIgVcNZYlkl6UUTnAIwEZ6T6Zuo9T3MSloAPcVwmqbN+JGth
WUhCq5JeNJ4wmGvIkvqTiSvFuEQhd+1NQyni3KOzTP8NxCO7cewpR4hQM/RWkLVKzMWc6SDCWZrU
eeUxH+M3+CnuyI/qBi1IsCmznoOMeDSklg1RASfGz8kyvsd3r8vp4dRa4OoOIauUYVUevv3L96pf
e9LE9QAWnO12ZbyDTHFBOrJwNaompIWUSKZp5Fu+AhmMYaBoxH7eiH4JloaNmaAJFskhXULivycx
I3b3mZYzTAHZ17JQSkgw1q5vNkkhgvGqeg7wbRd+DMHnYY7nZCRPRjhaye4OHMHBjDKIc5ayTuWR
zDe5q+Uz48hzFmlnhRZYiMDLJglLi7KXd5YiBDaK6IcK/gElP6eRRkmGWMdQp/9O/wjbxm4yfdZ3
wpfpfIEyk2UVNZQo+67n9UKJ08BIPqHnP2Ka/ZLSY8FwTcUNpkHaJTAxrIDV29j4gfUGInLZxXjK
iSot3O0r/UStmhQt8cHKOn30iH/smQvYBFb6yxcqVtlQCg2Zsb8qp4y/XR1vPCTWRo7kYDSt7ZFE
OJeYhoMmgb90YT9ElOf2r8ujRL8G1n5KsP+o133s8DDx+3t1Zv+PJfMlIiYNmF8znynjbC89uUFl
WX8YOs0o8NXUNT9xWF/tj1LO5Lh3uKMHK2C/QXKNIkdVtW6+kfwig5APpZZhbOmDakz94N0541Ma
99MmGkcU0JY7eCCmJMMAHE4dtOeFnF0P5hTDJTClYimupQHIW5RQ4KBclMWy2U7fA2y4jPi7rNf/
oMFYeAyF6bg5sEugr+tJwqVenaL5LLEl7zzCZ5tXVajbFpqmQb4TGtqjxMjBW9S4MxZuIEmaaw50
RMIoghJHRwaINgptCeOoSs3E7u6AnPhaVsb+u/5tY6QayOtVRE1HYcYe/ktN0QD7pzVHLUyhGfVv
RSXzcegMFbiRogrJTVfhBK5B2cbo+NUQEafZHQ73cB2sSONAhGlNMNjRVd9YYrySxP/xEelDN9no
iIkcvYx+Elp8iyW3YZ+xvUqxPepNPRYVHxLo5FPWc9yXgkaSj2UWSt4n5JwD8xWoziyvTqcWCZLr
pMUsW09r3jERm8KzNqeI5bph9AvYmtam3UAJ9ipChxG6TZwmXN2f2IFKxx+0k3htKSK5GW18rdO8
e/rk2nSxdvvPEIAWfZs9mp8GZoq6lmmGxD8whpHzELLCJHQPaRZlBeb4ypvzwn7Rk7CMYBgArtJp
zRhpTDxHcJIA+c2z/3+/ffBM/rESqRSqYBScIUyu+xE2hRKIxQ2f5Nh2zr4NS3lX9nU7tDji6haO
q2TW1QdpEHSFk4kPBh+lVAhFqAXMyd/lbtteowVqMEG7FZYCOZFeGU2EZQ3BVKGqjeU1qezs6BXV
bAgUssWfTWKORwqYjkHR6x9w8wNxVFuHe3u/tJOVMjafD9+mibnxibqhFQEzhchgayq+nomA5+GM
oqCrEBpjsorqgBUZ+Q6hxsRXIhb5CCzwSVys5Q/lUSt2LlcGex/jxiCciQxsGW6q5zDFeG7KJaoZ
V6fY0p+51voPlCJZUfozPkxnipJDLFZsEz5hl8VjlgsjICMIcJMZ7uxr5LtRz6hNR9Q7Bly9wCUU
B3NIFyyRZVg5rnekfpJgV3zHggr5IUS9KiERWh27l1PtHBv7Q5TaiLu3JIu054Zar9U6V05rLO/J
aW/XPjtIWDMps1PAIkjh5ahXM47pSD3FbXklZVKynSBETMpW3mIrKGR4DYaSRZ8A4cLusYRyoXry
A5Hq5XNV4RVBzqBPuA4fDK+BnrH5tVggqDiaHAf0Y1od19G45jlsyk0vFDS4OT9T6V91S5pS+FUN
+BWc2AE5Th24gdJvhHMVejb/izGXvTr2j4hiLbvxPKkZpaJLIwG2kTBXlJHIAufaQQummLjHAoQk
NBV8wheYXsyJMVsnnoRbiG/XucOYy/NUDpRjE47BafQo0TCxbbMp/RymaUxoFt88hlh/Y+F5Oex5
96sgvObvf0kNvjgnym9wetWojRZDtfvMiBjvvUwe86gpHpYTSGd4J2+6WZOYEHVeMVi4FHzwmy0B
EGeY4GDV6c4PbArMgz7SUYDgHhO2AXaRL+Evyz6lfDLKiSC4DN5QdsfLLCb5wey0yT2ZMGoLV8eG
gfxFGqwWyHmMA8vgJOhy3zZ4KlewGN0sDueXT/adnsv/2cvDfVyTLPTB72NQe8w+46a4tkJgx0Sr
/a8rRQ8EKYPDvS5iIh2wBHj8hjNadi40dXxMOa3CmKEKeIAPNPQbCUjDfE+Y8ueXkIcilGJrPmTJ
1Jc36jGmQoFYj1Ufz6RFV6/4DbwTzU9sCEC7tQHm/1/m9UbF5xYkStrmexKgLJZvsaOW6Y3HchPH
DglyVoqz5UldMiDBKS/gUEmygmUwgzHHBJp6jjyrL1I1bEv1HlEbsKC0aZi9KnS2r3TjMcOd8iaE
vXnOiRg0P5/yDIdxnL+Sb6xJHOyKHTAAKnY52+RPEeyMuXbKG0nxWJolSRz/DkSdoQT56aMuXA67
VkfI3Aly6YVpdcMMes+T4MpEw8Wa0Vl/CLBMQtZkdEw+oTdhxbovdnQ6Xfzg1JrqWuu3mipossfw
X6C6w3AqAhyjqedsqefMQudJFcjdqAWaX3lIivmEAYqW9QOw0jkGB8IK0YRlN3OdXdCrIR5NlELN
wpzRxcOw55bLE3ic+yiM53M2YPICHiSVfREenOkpljrFenT2YYgLekMUrN/54zOxOoUdN89olGNE
45yNjR1n2X2v2wvYc+ilt213qtp/dMWzCrB93aKl+rvU90PeNoEjrfOLvsEDr2NrUXPPws5lN2g1
QOV5XKeydY0Cf18CDggur8WMrDrno+YZeBlt1WISWeYfmX7IiigmxV9iL7EM9pEqg9juVx7dFYJW
BcufZgXS9zv+mzqMWs6vpa8Uid8PF03sxwfsWqaZbvpZYHhofVA8479sIml+whcW9jRWU6riF8ri
onzl87IW06Nxe6eoWdsVw1Qjds4u23qa2dIb2+hOfkwBSMwWGy76W9dv+fEG+fxMDyZhksS6sWJb
xJNtvRqZzJm9WhTwG7JRo0mk5HEan4hqaLeCJLJS7Sv5Rt1pTVaWwHqzlO37S6WY9KL/FAg7z1Tw
IOhkG/pYuyzzmuav8J7w2BFcMDXsFlW3etkZhBKvjnfwzzwn2veBn30UDhBRkJWBVPiBG05EURsC
zwCH0A+ofDLn1geEQMrT45Kee2+J1fZK51WlEwGHNg3pYuFlZMzmaydkmWxyY5lcxo7sqVf0+9aO
0vsq+BFXriuegLyP+3BZmGDPmVt/YVfGG0gmTHcEonVTbYcRwAHZ3voAqLIOfOMooH/XvoOU0AYz
I56X4qewetDShxTcQk7IQ8ed9TIwOtVW8YmmqmEf5H3qIXg1jW6brEcmPfGHbcRxz+vtdOvv+3gM
tZdP+yivJklCfpJJxl3kngLzC1MtRQUyhHbojxfpRovhcWvrwNWgpt7BFfOFAQ4RsjQRuIBW0aoF
ZRV7h+9dPtlrv+CiONDtU84jHWWsCyDUc+RMUQmGO5xfMm4qafKDxrJtqD+SCumd5gjTVMb4OrNO
qGnSs5POyytpQLTW4DKN1Yg1/mu9sFWw9w8qHEniCdm211taGM0khN0HRrO81Tb/R3hXBMJTe/9a
hpwpOuHJBYUkyx+6ibXcvn4SnIk4JAQdvVgfOUWG73CaXT6Rmr4oqMuVWoBw6Zu3n/a4Jfw9p9W8
IKQLZPYSPn5Dov3qCFHiN1mZ8WL/6vUA8Qj36DsejDlx5GNKV5DFNxGHK2N+cORRDVXo4FTTlmUb
ydutQsFU0bo2FsfQtzqeDfYLnTzLO9yg0PNxsnpo5auok8qnn1TtJ5PZyLRXqcdI0gOaR2W2EwN3
t7TcJquPsB2qwFTGZM36o6oQ2W90drVrg+q1xVkMtv4xwc848sya/X7sqNnjGL4nQH/jVN85Fbve
iJdBJe5HgxuQpJrpMUDAkuFy9JWJWRQYglEur8XOb4gsTZ1Ycdjn/F7bgGaVBMDKdZD3hXJpR0lC
VZEgo8xfROwjIWoJZH/dzehFcfz3DuCyjUolJJzvdCJGI2vV0NHrampXXC9mxGnDDQvGnLyyoJ2B
tmvATztDIg0Myl2c8tV5K93ZkeDgwZPkhOXEZnlA+Qh/zL/mcoxXP00SUL3TA2DUClKELrx1AegC
pN7Av3/CT8zKrK2AcJCcPyqDBUKI+1Ix2ToSal2Y0URb07y+bhdpNJTfG6tSHAH3L8HVgOruOjww
zaTJuAMIvJhmzAbnFShTjZ4C+oMPzmdw4RE9XWpKCj0rHbcM2QdIFHSnSXeWZpF0OgbD760/jsKx
en4gkjax2hGHPGW4Nb8HI2hU/SqBf3Skq0v+YcJ5rEhgq0QbUtUYITcR6CUZv7T6GwG1kYr9DunI
hFkvRTcOlZAP3YCGZCmRTYnrSyxLTcVP0GLUFZVrOg91c7W/lDx383ZXO7ZW7RPEPX9P/oh4bR3C
G7wiiLqYxYg6VxiaSre5FozTslp7eLaydMA9XFs4U0jZq7wRKHU7LCHQQjh1T5kq3SvwV8Rilxn0
hxRQDeQncMRWb9XJOg9PoYKZK2bY/p5Rm+yu1RPuE0ctkUYgAvRydFu5xe41XE3q/swSkKnfGbrc
kWgn+MqoEv3LOXvcGG702srfxgSCYucN7vGMHBKu+EOqhP40ipP4cgx8I1Xs5ptpPXddSu36BGyi
+lT77iXzmxFJYKHyph3EDeko2ov6WWHCylESNxM+07LgGbGI84p6lw9WuGwGJH1YLQGDb8olJsrm
o6giG3zHj/fX0kDyBVTGdzAdbUbE7EOI55HBg4/eB1dba+Pjqe2okNzDtQZstGkAzjQCWUEoM4im
tk9FBvXbtLEsrgVsaoigejWbFLA19aMdK5OKcMFNAf1JjFeoxj1O2q4/E/Hg3XowCPhksz4+p59c
zqapf5lfKZdHAXPy4jbINdeiZLqZGTMdA/zVuL2YjyBAS31FHsHeI4jXIsBcXBGJUsIgTQOtvXPX
m4U725+NyNVVpspqO/egBK4Ohw5v1UP+X3zkLzlmFowc2MkT2/OqyiNxC8qEaY1vIFe8rUqMZNSD
r+Tf8zY4uppdLPk6f+CtNmAaPNOTNyevsR9zDJocXv1DLydKgITPrN3g4vcviKReO2B7ekywfTYs
HzF5GlBlMJ+xAntaJvRVw8GPc/I0D3A9jFEVl23I/QmJepSvlsGq0Ggd4S3zNAduVT+cCIORgsUw
RD+w5tG7aV4kyFMZ4ySUIS9eDdHgPMoFxwJijlgekvcK3fWp5cwHW9p5OZDp7SqjLIgdVcIwz+/m
v+RmtyBP3Y599CfOaTocW5Rzy0X1m8vVQ4jmOWQtS5Z160PWJ5HsfVXgbN2UjDIXlf7wakVHlfbG
sJymR0bPF1vwgmxMqUSSH4k3a8qUdof9CzxwQGCkumxBizsSvfWr9D1ThHazdg/Aktspo8+6QEcI
k9O0DMGOao14KOUfMruLocn/MdVC2kWN7kp+Nj4i/MGzU01W1Fxz8hp9BYSUlTkDdfz6SYMAM0ir
vhCQEfE72VYOGMHJgnD1+0qAVV17tOHRkjF0iS5lPl8zLrgMIDAkZhcjlR2iBByqvktzU3etXzeT
r0c4MzP24gQAFTCaurEg9PgBEBkF5aUYwEIB9FzIlkhGxL/dtOmoPofvRfFLXbmK/criEVGobaiB
JHY/67cxpxj+uVytyCBt1KOEdhrBRgzw91fQo5NCs1EZOB4isDeJw/w9h3EhCcoWL6dyMepdUbJR
E2YZaveLgr9ZOI3sOgwWQMB5RkvmXQvxzB7xVnMv03AFVKpNLoCySqxdHVUy2K40w6i1nK16Hmfx
CmASIFrPBKhoTYVVss+m9A36zGuN9Ky2/MWjhtSr1pGhrKIY7b+5jJmI+EmDjykFXX//XLgTI9nr
ofJ4UI/b3e2Q4F6bHtfddhxthNbL7u33SBrPRsIF5tO7XoYBtzqmzE+DDTxW812pGQbA9qcp1l+d
IvIGJ/2mzRGKQj7DTlr9bUyf5AaYbA5T1u62+qjkeyhj7a+/TgRAqujHdgehN9R6b5sef4djg3uP
Q49IU1c1Qlqlgie12//oZMk88w6SfiirajgLhq9fmsXOofTS94GN7dbVktqNYkIYVnkVA6C6AQqE
ugcCtAgU0411xBEbR/oDkIBYtQKOnuTdT4nc0PdNfHA+T/W+quIZf3iQeZjJpa34VzMMjK3Baiqh
CcQYrxBGvEfQ3e+q4CVyVG23r/JmC5+kHXbKVWRRdSXGngpAiJoUd1/lRptUK27HlWUD487jR3HR
BTJtLUsc2wjgRkHkC45n0Q9jvQhgeW3Aa8VeSydCWBJ8EJAeLbY4zNOWt6E+e7P9Zp3bzcrGyr7p
lxexdIzgsEmcHjhT7OchZ8kTpxj+3Ceu5iPSKa8BJTjaPViS4OYP5MljCFkIkVgU6EJei9A3k+5Q
1C8Vsatc3fK4KJkE1JL8JJ5mOLYNCrC7U5H4S/jcPyEQM8Ws6DJ/8W5kXoxLa4lhL8s+ZjerFAin
sKXdnrcCrFcl0Ox7wCvDeYrYi0F86Kx1MlMBgsHjjoDSpNrwaPMwLe9a5XE+Q3GqJpCda8brIWj1
7H/IplShsAwOO7z/mN8MC0JUxtWb4myP0J6T2p30akghD860+5Jyb9fNx12qVVjCCDShFLsEZ7+b
Dq07PUV9xLGHsdejCRYt3JjXZPSvbzg1MsbUea1f/0hF/7cB2aTpuWcWpRmiX8qqHiTzN5MfBg7E
oURYyUXpodKjbBncBDzNwJw+iM1BQqC712nFgnaXdiMU8Us5fN5FZMIeRG76+/Osd4WeAPUeQJUY
1oq4KKfdCE7hV7NBz//akZ1CSGq/MOTjYYYqLOTwkJ3TtGVoFcAkfZBIUQdRDTotD+N8INs+M7zO
VJj3JNo8t6/ORZ5vRWgRczaLM9JKZ/+bBZRbz5MVEg1lbFgamDT4tGyQx4409qm+BRJyzqpNT542
pFiI3m9XsaJchmdBouxTyEzJsRntUqW1v8TJEn1i7439k+OWNLCdC8myOUcJam7nYS+Wt5hAFWD2
VZDLrKxfMv64Ab9Wm6EQ5gMTc1OeeiMPp9+Z6D8n5NGkv2Z5HmmMSWcSyoAvEo20T02kCZcvd9NC
3zWtJL8sOkSbZbWUZnnc2C+W7KrlrQH9gDm/AShdXfver9fb9iAq/yS1AWCTo55ajfBZA9f0jGQS
3SNV6YuWGo2EHzqpo946/zyNS3HyF0jkv+SV+PX6Z8/KB+rSyrlZkevIpHY0GF0C8xhra7XD22YL
QyQjLRKVnuWBExpUkaoKDLjdig2H0fRq6abTh0n+eVgrsZ9Kb+hgQ9w/YiPyszS65PXJF0O41JAR
oPLE69sNl8L3nprWZ9g5alaMsYFg0E6QwVq4yeKK8W9hvzJJ00Jc6QIvqndykru23K/gCafP2CwW
9mj0qmjmyV4bYL/ePzRvIwTk9ObkxQsCt/5Ruq0W0kjYtMsslawNH8KSq3FfdFS5S4D11VzN4QpN
U27p3OcS/G1mFwPsd0PHtlwWIJpyZbPPatQewLZNH2NIy+/QTkrIN6q4zkKuYBf5WypH2TpdpLb7
3tt7ksC8iF6r2eDPsTqV3vjkp4ivPSS+rtSnCDJ5N5PWOctDpNLLIkRxm1+XnYQo/iXfHYVmS9vd
Ncehy0/UfMHdC8jWrl9YVOv7IVGq+f6Zelkbr/gwe4XROtiXFX1EH3iV7rUXIL2KIu8L+jLRzVCh
k6wbwoG1DuqLjM94vhjerx2d0Qw5B/txcbODEcqQYxqW7+kmeGni2ju/Wi4x2lb6l0gY1NZuOj7j
lGu2cVpn2nGWwVOJh+ylvUt72OPPg81Juj8n67VesmXtSx3hGFlLdQ70DCUBhMnUSlxw60KPR5vM
5GI+5iX7/uRZ/HSXLT4YBJPX6HVSJSyuxTxDo3uOYbCPAhSLl2OWEoFQiHXyA0G6yhyfPMcDR62p
bhr7TypG7tsS0pjg+K+7gONT31IGb5zuA1hgt/3rfInJQu67c/3/9gt8zoYqw8PMPL8YDDKssEb2
xD34J5B6Iq2niwCeOqjqqsegMBIyDNL51AmaIEckLz9YvF2r2n+DkSRtyk8ky/zNIhi7ApSijH47
QhF0w5LmPaLdsAgjMLqGFHsBKnVBLtEtfGNJYPrqdZ35fF3oKG5mU5aydG62PlhSf6BQhF+KYba+
plqA4XQLyhFwm4yHDBY5rzek6bZazMemYgQm0IdeCnl/RUcSTrENHxiDW45W2uX3C3ztacbgKfN6
BJA4DE8VspfPp4NrYqq69urpBr9jYZdawoe9jJ72QoGrpClKleif44ojt9GeajpdtVrkCc4UmJjV
sotTQSgNKKk4tYqIf/fApK17Y+RzRZtn6LPmz427anIvdErqVqsCmFpR8ek2wDi4fG5gDIeVkdfQ
wD9+5eVMdmZGw8CWJWKIq8S+JtkN0zb1B2kAJDGDBPiJo+j6T5MnA+y50lp12bBTHIeLy1B8fNQc
5cmv2sIF0XfVyfhV7zxU/aWF1Ps2EwvmycJn1Kb1ThPBfblk/4xU00C1Fo0ukaGyRqDhBC5Qyd5x
hfuiFholIFmSgN4Ep7llJ8dR1j4/BsY+Xko/3mrLQMifvqKrDROJqa6ec7q8qCMMLCAm1gjvS+vt
EJlkHBflNd97WeXb2u0SSjo0VOookV1QLL17kpL6JnNCh6jvm6e2CoHg1TY/HqPXmM/FpgLGWBCS
6NkJEtPZl6i8IxEUEHMbTYSZvFDITbKdrBCi5R6ra4Y/p8iKRR2n1uSa9krl3OXKMFZ7jXCs0J7T
NMk2NIT8ldiKFML1tNQ0vpZ8IxlZMVvGkoGtQKW3Px79RvSAyx3cI9C10QK9LTirWODUZzQtfI3B
szY/04SH3BQPUW6WEoCMiY+mCDfnHcU15OuyBL2KJeMSR7d3xzfIPynRajbmz9jzvT/ber++ShIA
uEsKXvEo3BRRZQ6q1sMDxniPfKjXgHhV5kg9Y9282y4y9eqIqVox1Kk/reDgnLBy/zaAE+1N+kuk
it9G1gBzz1wZY6QEVQ2bllKbpPMCz2iDgRHqGOcovPsMWnmaetx63UevvR535Ebsiko0sDCf8UM7
cvMp+wwm6lCdlA8S60bQfaoG0G4Bp32xJYCvc6TpydecGqBY2lNI7avP8Xf7uJe1X5Q2t1Xx4iFD
YxO7xQKcdzMcydERaq+EG7k8XjL1Tzus9J7RQWRQdUgXaEK+loso/mj362yksSDfNgFyp5+yvZ6F
odMIf/Ie3D2QMIGgP+UxuRDAi6Lkw+vqBOjXA1TMQRguu3k57L006mE7wAOZwjnLhcONErREUuBi
GHDPsG41GXZIBC1Wqjn9i18dFxzmr+zEHJEB9LcDjdcjtWrfv726Ur5JIV/pj2PzprPIAZNtgJcu
1O2IdJgGx+MtYunthLXX9BT4jD5jza7nQ6Z+e0UCsrUENnDNnJdB+4mLdadPhfHlMx8i5QbuXipE
kQ5PMohjA9K2rhEHaOCtdlDmEzULW+3xIj0g5vFyAUtCoGXO/aVzNDynkhg6irmn/zfKY/zdnpkP
7iuOT4ddW21w+cpHDPYA5kDUAKV2CouXXbx7sJxKBXK3Xu1qWNRQttsBU0KYmx6cjHjr+FfXimNr
vvAJwSpdietsnE8Bx8Qnlc0vAwPMmBRpIoyU6l5/BghpzRUnXYw06VYFd9aAHnDEI1xy5SfNhHRo
h5MmqZcBWZmkEnrYYrKPsR8Wwuoe7v4VYA6rst63oAgEb3LZLZ8NTYc1N4PS+C2LfGATVP2gQydM
G3ppcARirjfKEPwgXgLOXsK2g8gHvLcbwhim5XLns8ibU5D2yWl4AfkOlzGGDckxXN0YV4+z9GxP
Mkkle7tostdidLcxxiTCOBKPfacldFWfnSV7SjiJpnQYTso6kSH/bfjnPVdh1hZThOwyMrrnHnqa
8OPP0yrgDtE8yhgR+KzX3Mygbl5A295K0doUC0soySSvpRVjd1FjEMTIbbRb8T73kuPkVG+HsRkG
VmZ3ElqEzPu+ECm4aX4gdAy71csHji5LM8BvgWYQCpfzdvftFhy3BOOz0BjbB1sZbvmnV/mOPplN
j2Nhbxt1u75Xyix7pvbpCIVTQGq0E6GGQ8EK8cBejrkanVBoRlnOVoqefmyheRQClHrqk+WCmTw8
VBTezCHSoKOj/LV5rwQNNCA3ZYVj1s45qRtnMI3j/bAY5DQAYVSbDa8smCJv0qa3c0iB4MSPda1v
XdaBdU9Rxo4NbQC2Cs6Q6M52pxTFRnP4its8SGxLK9hzfs6UW11iMQA5nNdYHo51Nlu5A7pJ8ztp
HRsqzXzx+tHEGvloMoCR1RhzTpf1rhwf61bOTFLSONL+zcgPLFf5sLLHS6+cM3a8+G0YFv120tZN
Ghz8LvYYrmoi/cA0v66pcCEvWKiPDAJVTjs48s21351CYZ/YvVSScF595z7vZ1CyTLv/4URAaVq3
87f6FyZUuBzuECdN9jJvilKzz0/Kz8Q74A7CvYJqBFZXdHXpi5Uc/dhEfkIhmiAgJ/BGIuhWeBZD
5xPeCNPWLiedTYxgKajgW9PwVNvAczXGWhch6hleV+ctXxOQLXXT4HRDa6AbUJU1b1aFzZJGnYdg
cgWGyEI+l1q5BnZ/IGrHI0Zp2Eq1vq8f+b6JvzVG0x65mMWD1/AWlWNAs2ZjhTbDZ3nkHacEFo3H
O/s/Hyt4S/Sht10R89M0QP1nqW7g1A7zzrXVx7HPt257Cl+OmWK+1fI+/iLWG/VQHjea4HE/aOBp
84wC9FhBLrgQ7OrxD8rZVXcyFL9m+qTp9eXwc71M00zA7+HYjRasOpvIGWYyzQfueOlBUhFxURYa
9Obpzd8lxy5xwljF/rKZZPKhKOn/SNI6dkfxuNCWOwhAVmaSKU1hRc8w70Ka6iQmGjsz4AjxMgXS
LrrOkpFzUnGKfhy3tRSO7MomNdpiVL0pseBV50s2UVjan8NNLXzKnbkh55t0vT3+9A3WEWpMD/z6
+eYzLn2t0/x32AgplB9UitprYUBI1FW7HFuxf/XvurgcaAIz639d2OFXgESYg7U4lYT6tOcgxUWf
7PAPbbeJmrss1XiA2GrikKzfdjZoYyxK1uRs83q2CqE7N+bmSCqGWReOezI+WXeh1W9NID4+/bEP
MulxCmHBvoXCUalW+tv91rJYTFez7O+u6Qm/0GK40GjQ/rJrpg4kWOFv4GdIHrh7cffJVAS2yjdP
mtQXPshD8EKz9By8ar9LLyJNevUFko/3BVZi65G3P/MAjQG5Tav04eSnHBMa5L/4uJCxwYOAaWn1
lOXo1XohWicqSa42P50JVjCSKVWJgyKfD+q9xI8RDO9MkNhTB1b7vjeNY89ltat2VYSdYiqUXCE2
G231GpBDhhH/tl6askOJ5QEwKUIyittQIYCbAI6FW1anTNr+i1Wh4ei1gVYlYUSqANXcM/cfxKmU
rXGI5wZ9uKER8ZnAbWcGUFx9LUXUcxH6YGWzIMJEAmrYYGol/aeIOz42Y0UsnIlDVnoIfXroNBVF
zyNr85NKJ6yOnpCzJW+d9nLUW28Hqf/egJ159DAKkNWIDGl9dBOsV1BrMSGWWpzZs8bR0yVeqd4+
biNDRbaGvMkOhavMY9piUulhJWqHaQQybhHLIM3dy78cSsA8292a6mX3uUhOeeCZVG1JkY2scS+U
vZSixnzqijAiZMrB5Y/A8rU5nblICFATzyNAVi3c2SsIy5FHnm9A2cCgVqRZ0UXyGWMtFgpDLnvQ
i1JiUHvvKISCupSUNDFSGhvnSw2mUfWQHnZCyCfyUAloTSJ+oA82FWtZKdoU/qJyzGGgoQ755NoY
dbXFsuEOX5H5ez5EEMmwc1tz8sfBJOQ/Bd+b7rOF1qhL7IwFU/i0wvulaJlP002LSmOTnbFPsSV1
HFRZfeLzUeN38NuR3fppCvRfd0F6V1tx0Vtmkfbpt4kL1ZFUts0JsVFDyWOT7N3ZfR3U/tKExLIE
n25Sa6fK8o0a3gMTdWVPnYyZkXTm3j7UvyKszqnAlJ04wREp4bIm8Uy+wAE4euhQHkI7UPT1Rpfs
HRuVoIWEagsVDy8r6xo8ZljZELndUPHKD9klVC3Q3rciXeXzqIzYfQq+g+Zfg1D5u7VtROkug1Hk
n6SRa28c+JlZ8u28WnTcPz8dVHwiS/H9U5vfg3roVet5xWnz0RsXP2HSkGg6TCbgqnRS3/sh31sm
FArMCbR/VMGHUyUnaxAamHoTxFFHMqcLvyAwP00Kk0UjrTfns4T9Bac7p6vCLowQconUd+1V61/h
97TOYhKbT+5tKiCp00xJyYG2OdMrZQzkmzG58iI8Pq1HaPTmh1Oy7AEgs+/oLb/d4nET4BHFD9q8
7n7/HBVUA49IuO43QvbTyQNB/a1uiqmSsBxDV57DtLgxgpcyGlicGwZUfoBX+mDun4lFSwdS0bPG
IVVZj/YOw/367jwc3CR63CvKNXd1MCHgH8ET7ciWFAOyWrL9jigiZn227BnhY/DTxIcgX3UeyHpQ
8FRuy1xjtYQatr7HE9NdaGcVmaWOA12blFSJuuZ+yaR+ti9kp335pX+haYnKy73ki7i1w+h1EF0/
VXq5L5tdNOw3BaN+e7QmyUCqjonA+QYQ/H9AAc34a8Ki71bCAcgEAyU44QB0sVfbFE7asllSwtF1
1JxU6CWCIT4viub0tkPvs/m8LNLmZsdhLMtloZbPACv5ySxBu/8XvyyQlAMpHU0tJEyeXzlMgMuk
TPnfBifKz01LVq29tjgICbgmE7CwwAiCKSz/3P37+DUav5O9PHsG9bWByNbX3e+yNuANpYqje81M
7QC64ak1h6P2NiFogAe76R8hhsDKxJ/YwjQDlDMjYsKuqMs6qSlOEilW9VYIU3/TwPiVTYca8zTd
yyokuV1UIqFSBF4clP3f1vpnmrK4wR7uthtv2ooWCycJlb5rQPjqDQ75gEUqWe2N8oQ0nIo9VkQv
3iF/FcWyIRfrnaGJ7Em7pgFCbzZkD4K3ro8iCILgmVAMuY12KGn/zghnU2UOVvq4/Z60txR9Cbve
QoETa6Fql5mnWOvgUUv98ZBeqMnIUWrvl3e+muXPn2cdHoTlX1NtgBzl8IklABa99EV5d78g2l1Q
b6CbrJAXbsTmIRmHpMS+HdmF2xyfyroYZ3P1fWyLrGWbKdtvM6/c6gLuTsk4rz1T4ngWFYytku+8
ZKyQjkwkSXnOPX9iWoqE/z6bM4nDc564qF2qoDaegQCNeLgi75eHH+MkpIIOtzKMUmlXy3+Hq2iL
hFBZl/l61xtq2LXEIRPXwwcgsSP4pQ+TFy8GvSR6LhfMm5AbtPP0gMbeNEsPMUI/EDMUo9ETPfaP
0FWRrjQ9bzI6euFWCS7RQaLTgBXy70cQplcVT0sBLpfKXCpP7WH04ZDFLkv5w7RZT4IbIZxycitH
pRGtBJ/L+VcwX+dfTwJ27jxg9cdHj0TRMlgiLRpl0VmQdnhbX+CKK4N5unmyr1mGlcw+OQgeFWsi
mkZ0StFUkLM39vg538bUFqPz7190mF9m41u4kTUtnmWtjguym6XR5WU70SNOo21AVXDYKt3rgY0H
UoM1JQsGD3QU4j+jcPgny9WoUcKVTT9fvAeUF6vg1q+Hh4TY2AJDEvAKMjf2nf1hOgj4K9velLW/
C/oNgLI7xkX1qRJ5GDPg3tdHxSrchqjGgQDgUg1d7M0TRKyJxWjYZVBAtiH15eSvZ1waPrEe6TFt
VlKJj72cbf5pC5gsZz4y6pV49Fb9lyzcnZLz2dEb5vWJLOf0L4fZuxHcDpSPXmZpRwUHGRbyvo3N
/YoPRQCJv0nvspvh6Iqsz+erpMpU6lD2HHq16UV87+4z+1cBRSUoVH9jurTiqPjpVoPKTm6JPQu/
pvxKTiS5P1BSV09o7J5Pun//2Bae4BFR9qxzzx1mfN5fCuAqS3zo69n2INaWCRDy7HJhLxAUTMP4
0Urzlljg9jNogV7rNpQhRWCUjHBqkcwyqYL0L+HcNK75j08tVR9da46clu34DXByJl+4Up/TCGtg
DTTXqVwFK82pUMs9dd0Wml8yDkZvyV+hNnArhWHulJ5Fx6CRhrC45rtz4A2FoUXatHtOogIYBPQb
xO9RjxIr5oVyi3GsLy0N4RuF5IEVpiZ0JkVZPrxOJPjQ8UtcN51xuhVnc0by+vHn9DOU9NKSWKdP
rjiS/hUmF1M3MvyGktd0AFkwwGUdEggKkCNOxlNsMTpDkItUzRdf3Wd1PcoZvqY1yy8NcOge48RY
Ot6iTiOizRLqrrnNc0V81jEgO+P7PMA/bJVQQBsjBo5lbaQes7upyG0OIZbLj6qm83JXBxtHg9eD
aNy+uINPBWKRwkCxiqALxpb40o8lLky/FeYir5Orc/aC96MBVTJmXeULtnb6/hm1ciuja/5VwP0f
AwZzqGmhif1vFj6OkZRszSnAeWiQrLjoMj9erkXcpdAZ4EQP26h8lXcWPjtJJVINbGnz/rcxaLFp
CbsHW+onzeRKK3vOuEi7IgcQrsTEPaS5lWBGNBNqvpeI/a42cTjesw/wQdqACoCcfeNqO3uBBoA5
hTe2U817WkCov9w8WVymd53qSCHL/Vd84CaQbT8iB1Kxskhv8O+6YFOFxc7rKmGGzrHHvno/y6Q9
U2HsE9xUgl8DRJ+TgJh13nDAdrTpbAIjJTQ1HfXctizIZ5XzjCmRyDsL23J24JaC4tXtCSMcOY2x
/6VPrvDrgJ3NMyzk5v/cfb3B9fstE4ke/CH8hNOLQ2ShS2uX/jOB1JJ0gwYpStXt6DUomDf29mtA
xlVHsLKkhserivGW6ajuch2yw4ZqOuAsqyzl01Hs1XXHkpwa4yeu5D/J1ql6EGgRR0Ibri9s5Wb7
aDXVvz8Jt/zkTd3GY2G1AAyYjzbA63hxorbot3Eu8mmXYP8aqHsyqDLN/TZWgHOoTZKIVNXrwxIA
60EAq5xKsWBDWNyuneMfVp2LLfYUwAkgF14b+07WiFfyQ5zlDHw2WQvTvv6bxC8jA3QQhtLdDolB
J0SCHVO5fGGRw85IjWeA2GptfxzPkO68cgcWusndW39nlVk1Tm3d5iO77iKAaCRd2gJB8YD6TI4U
ceRsBwidCknj7vPB2/7W3NrBV42y+CoI3u252Z/W115Mi5/h0CIgX2834/wTDKeNO+Ea84h+wLGb
yKx/YEz0O7wlTOKgAqS08rehweOJhUPWmRJhymYCtes3qcxP4EOn2ssWZUFYxtn0VUZ7m2DF0dq1
sRMfbEqD3Ce6G0D6uW01gt6hoNrdGhUW0M5x5dV/2TR340TTUO4boAR5iuPVTlBbOEKBx18CsKCF
MCDDWSYj4yGnRzKPwqlfFxBLo64hUA99XXxwDPGJthcvF/Gs6xWnY8sY+ICuEsZG9A7ncGjeBgXf
IJ0i/a50qSH0DELiYHLPYp38hCvU+045IBTe6EZ0cQcXGB9SxXNYGLP6WvOAztsPnjsNn3UnX9n3
GJKN0BeyN4ZCuq324DXJ+713nJCSoTlubcHvXKn4Ve/6Nz5SaWsbQFzoJX+UGRnMOoL9ufrqveo8
4M0sbivrEvIcLy5sV8HuEH/5NVf28hyfNyM01R7anrBKe7JNfbw6MJz2FH/AUviAZKKvutku+HSt
i91XvbmoB+2RD+cJ6SWcq2VWv/8nEwCZYXr8TCnKt9Dsb8L2dvG89V5KQRwwahz0Q/3akN+0ha1K
eHjQntULxNco2FkWxXwMr0dyMwA2j8oaRikiiOi5K50z69ldrNMtGqGiErY/HLIPciWCNWMzd7eg
yUW2XUR7R8ObQTsix+eaazw1SN4nas5XBk2JfkzHNTtnqZMdSkzNi/fgM54CB99Cf8j6GSX6Al78
fcIvNj9p/EDukRmJaMn9vxbqNOYjzTQYPMG7wq/79ii+L5ErtzoAik3/J0ZhrQ6cO8QXGbmRlVWa
jOq9hT1D6vAvW6st27Fa+Gvl/wDKgg86d4y8YhXKF92bab1LZbbqG7Iui54GM3Smf2SQQtWejZxg
xwwITTOAzJoUwsqXp48rQ+sXjbnCnS3KsYvFAogy++R65ThtVw6wKL3KrogEYAd+kd8YFXfaAG3G
aBYHeaZ5eMT6DZHw8euj9aYhlmZjav8UgUGZ8pxhRlSLJp9sVmWOax+jHjY6PhjbYYrCR2XPBK34
3wFnUucbJKwnKCk90K5u+NS2H4VT6/w5P73LgcrZMKEJvHUe4Vk4DCjepptalS97MQ+gSJ/AiIKh
ogd/051cav64yTbgwOxAVB+a32pau9ytrWRqxrkrrVLeliRahSUS2DXfL7jiOUXFy3BerIAA7pZn
n+w3F9Nk4V6ZUEiL5C9i5KGql+cTHg+e6oZVYmebEfGYKL3eifCMtDRSSZ2URffzKTGowidnMKcd
RuWM9ExAHLERlotMW3mVGo+7xvQ31WM+vO6CLcI7k0znftM5jR5KOmK62GaVbzUcMv98FyDpSBcS
0ofD5bOliEXfbZRuNHDU6/L86sGv0eC6TzgWrbPoIEJPWy2IKi7ZU1d5JfPrpgGcGr5ky8PxyheJ
oDbj8cWjPhGaH7rk/FmDr6USnCZdsmpJkfCpNmFfnxKzb41tKuga5J05mnSAJz12IVxDOC8m/FdG
ZBsH1XMurL+6Q2dwo3LAK2PCB22e+MRdMngkkO2QZiFMrOxw7apoFjAQ1wju0T9XTqSO4hlEa/+v
wqvlYRPArJ5I/ldUWf2eabG41tfM5/4O+JRm9LwKeiMHx2D8L1cPrNQSuKv3+2kdgKC7Zbnch26d
MyBvMRhOq4jzy6qRHBznY0HaPg8lxmCLMoazskEwd6JExmWp6LPwiisWObOl980YBVHThxI8az/J
w89bHUzgepXzKdO4M4ZhtBtx5k3earHYHWC6WhO1lJvol9H6GjvKOnvzE3I8enHakMHXYbwx53lr
4cVL4v1EVhpGlp3mOnHObw5PyY34BDNdturOuHinoV3cbDCEwDwmJ/VSsXy4CToqTmFDS+R+pfUE
6qnH20cjNd8cVKYVIf/2ksCZg9is71oDRvuj7KEMQCg7zH/pQc5tDKKqh4xx9Vkj0xkTPu267ioZ
G2yutEDt6RIB0D8aCYHy/AcFUBUEl5mfPQ59TkC0xQHsb4IGMGTuPB+fMIG+9Im2PnEKT3Cnrxq7
8KnjoGqULvch7rUCIGQCkMC0WwLBiYs3KtoE9SgKBadw50TWMYm8IIAF87qUMrsEHjA0+W18Lcq5
fjx9m3emUJRtQaJw1mSWWgoQfJpocrvSJPfMq8K8o+EQ1m3VQzFarh5MCQer/mAagqMiJMBTu3BD
0DYRg7kh/DowidQv9x/MfOnk/bRJg2AK6SVVT9rsfQDsIsSZLDUk31aQqZ6GbamXbmLobW4Zc91e
zWyM6Cmi9dHkEdARo32ClLJH7fle5y0M1hQ7mL37II6XabUVdD2p8vj+BiADz0maara1pCmCGx2y
BQzKMEWdSI0R9YM1XGwRW01wPOS3AFVyCVw3+E+5XuW3sE6VxIKCH0CbYqPQpJAK3Y81/5ob6ipL
kHJLY2RU9AE2xck87qY2AdXZareRzX/3KimhoD+M3+yVBcQqJQa6HXAKP9lZkXradxCaPoOe3eUz
2W3R5ai/+mGs6e9ogm6SQtXpGWeD3DApYeD/a5eFAehRC+PBnM32bUFc54S8IdpsZsocpyKh6jD3
mhxYJ7QKwo79DptWqAuDuw5c3sbDXtjq0s2f12bCsv3qVIuv2KRK3lqLx/eSglTN/hMmX4/zYWoN
Ns714bkL6iom2s4MJlQRspVx/LKiW2bmLYW2ji8i77qHWSkW4OfJm9ateTbzE8pO1s790VoKndWD
t2sXpljk4yhcp6OaeVQO21hG2Z0SbtE6AgudetWVsZt8+EviN4MNZiRGsj7NvtUaFl0Z39LLOW8W
c5TelG8b89I/kJ8RlZ+ydbUavRzEcva30jOhtviHGzSN7ID+uNdPYr8ktj0BmLV84Ulo4FOhpUEw
i2SH35ARQ1/artWR7CZuHr5yR7l+K7h/8SnXkTjf0MwJSQ7ODASbFPtVGmks/PybMBptuFHsEekQ
NbcySMyFzjS67x8+DTBI5DoY36mKSmCyXi8p1RsAvhAi7kyY2//p04b3Cx5R6vIFnLzpw+C4DgJJ
e48DIztUBz1yhcE7nhs9Kgk1LUuQaZh7ynPbeDrqHaCVOy/FcJJTH+Oe9bmcr14SAfkjoLKULVgk
StKeiqTPJzKCnNJGLckxvp4XNsB0KxXJB7r22N7krBn/0tobhDUBZaOAUieY4ARMI3OLnNvmQJXL
NhcKCwipdbKrSacfbJBZF+yISAK0kqHVklQHjI0=
`protect end_protected
