-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
edChwYygz+toEHq4VPFGfhaZNEsHEqabu/Otf5woyzhZkCtHKUKO6AXSufiiYlUq/G9sTTdEtPDE
+LrsatNjvfTGyEuJPNbd6vfxnEEq+Z3Hqbvdv1bRdOsYatiur7z7ZMPtCHpQ3HJ+XTroOS5y9ajc
dbGCSo/MMNpE5rlAVrwAsN4C4cUAAy5H1rD1e0se188Zb7pnWdPKwScLjPXbobHWvpCuWXn2L9MS
7TNp/oGsWYfD2+q9+vLMOqUDGSNl4EXWj3tqfmIbtPbUXVWBEsJ87x5zLL5y3SuZ3ExN3ME2jYLM
WYe8mZJeI1GOrpAuK+gmkyErK4r1TRk/Iu3C+g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18800)
`protect data_block
ixqLInXYI/poy2f5Z5/VgVBZFfX2dEOc07XtJKTRhA6G1ulfz4aEq2lebdZ3mfbpVpmLwNxUVei+
NkEwfTcCRvocoUVuXExb9C62nNDJGUFFWUwCV5788nf+8fDRXegA9uolQBvSCtv6ic9Jfk+FXB96
UP/R1OmFdCPn/dC3dXfP3D8aaonLD3myH0oDYM0rA64CUcg8YdLYGtHDH8k2aa4yTmJHeB6nwByV
uzD1p4EiDAaL1wCP7MCko1JObmb1GkHkvWYGHy5OZM3NiXglJcvyYaH2oRpJ2z/KwYiT+Yr7KQTN
bD1whZOX+YzEPd/Zu7cuTv6pSQfRGhgbHkDjKPRwAAcWXAt6jEjIt3NnKDx4XdJwhnh3Ipcd+0MN
yDjcDkxhwuR+ZuoZkmVKKqE/qCNw9hpTTpAlvG0Ne7zCwpNEurfQKPjHAPKPRBEDSjZqE09evKUg
R1wjd1E492DhyzIQKcy1XihRUyJzCQ/L7Q6qHhM47qMMqvM0H3nNFugxlx3hIL8CNuBgPqLNhOTj
4hg93wH+1MXNfGunaSJJVWKPip7FM4Gl/Qio135uQW3KnhzQ+bSthO8OblXvW5/6L40nG12yaA6z
Fn4HP34IQiWoFImt2f+quh+BoFNQ4oE9HzKM9/vO9vljcJcsfJnBA3N1PykH0qwATW9yL9cmw3C0
xRtjXdgxkaszl+S8kF/UXQ6uuTykZUleL134ggwUDIHup+KE7tbfdyCLXUJOuRyXCgDcOLkw/THI
B7eJJNkU4L6zU1M4ePV6Zox3Uzp6ljAsLxLbUNwz49swQS7hlV/l9Bp2Dj/SfswrMpTH7kdgMI+b
ilBKdY3/KqXZSxmWic9Q9Y0NEZ8aV2fWKIdniTl3B+2iiRnc3P2PG4cQzbhomFXXNibFQTkuQ0G0
hd8cNRv8cYEpTxUSV2RdoQolQJ3p67c6IQuDJiB41mgEFlPE9va1bNuQ5Mq7c4flHoPQHmg9pkzY
eLtmMSnxNgNT4r4DWIAnmphKbznPwv2Lw1ZlZoNC1JHpjOEwIVILogaJ0yord2o2+0rnCzHs3Mpz
lDhAtw6nkB1RKree7mOjcG1vtBqbelVyYj2TvS481Sq5IwseRkQfP+p/81KOzZR7AwAzga9pd6Cd
DstnLEmQ1GGX8Gq25Z1RQj8eLvFaICtjGbxoZxbOjUM7+uJVQDyGHzhK5OWRQoIzIBo2kDM1I7la
HV/LQsm+KSY0p0BVCY3bX2PDUozqs1uwzCzA/TtqxQWqJBZ9cZ2u9JXOldY8iTx2vcnt6sULiTco
EdgiTn/vsumVMsRHqyIwBJIHExxvv9dukd1T9m+vfaDYR5uUvTuSTSuu9xJ5/DmZx2Ma0fBjrApj
qB8+KlrbiXjeXc3Spo/h8Dh1lYyFGALXDX9+JvFuY6leOdeZeH7ktQ0NJyLD3Z2x1iU/Vg8+eDvU
Cq8KETHPbKc7sfhUPxOfq8Ohs8VTWjYAwL2/SXls/4vB0EsSqJpA1kkBWVs4aUKs8BxoArO1QVgl
YLbE41dM02SA4S2v+o7Xvkhdd6+Gf7coI+csuPOBk9pGO1sydl5a2fwhutevmGKi1H0DN19g6kF8
QZ5DL+qrfnCMYSJXZGo63YewPsZO3wKzk+IhokxI4NNuf36NdMTei1ONlRcrNgBMZBfwuEkf3jSz
8DnHmAfXO03+YPNB5VRHnDS14kIRn9jBGC5rOxCkeTRT5yjMHjKIiIvX3MHB691snCD8MwsEqANM
KCFCP1PL8MyHwaUr4Z5W9/mQuhrZhePJCqB/Gu8bIDjK4OaGQWbQ0al39vFi5dYe0L53Dg+W2OiE
Bxu+Gv4aLKIjxBCjKV4ZHKOOzzoVLSYEJWOsOiWQfVWs9jKiOyTolAIyH8N84LgUnDLyegnDumD5
c+PbrxY0pkcLJKEUV/tr4yfbLN5rRXLGarbR4vwBpbw/dURl1R6RLq57JFCw4av1JRby6iSXEBbl
pzCXn6+zvgSO3T5ILgX243MXp2qTQR00hAmlYLhfPPcm3jVztwnYEHRVblnIWDcN56DUjBPqTQfm
e1ssBSFXe5gQVSI1x2FV2lQvBu9FBMnlDV0wRIW75pzCqup/j32x72e59O5PI+Q1gIgMVWRo2o8w
TFQMSpDDgtUTzz93oOejJWLeDBe5S6mt1/OQvDlBadXNZKLI4KIZHQvbp9smYlxiUJmQj7doOx9y
H9VAgnBxQbf3KmLxb1fJ13YnGwDIxRtmUuvXiXVIsJxp7aI0qrF1/4vGRk5Inn2HUX3ACcO8+lB9
B6wCEc/jDpXnIzrvowdQ1wu7TbzaXqFDgDOdz7ETMmiOAzlOJJ6PYtCqYpMLwZgnJwMsAcr6gTlU
KtbAkKelHoXbGDBbiI4QinCifLa+Y2/3YHZ48uBpuJWD99qg1n9kNwZaauc6FqKvZ0eHGm0M0KgZ
PD38cne/SER3hBC3agOgZtPVFSJaaRwqjOT+zh4i+yCZSa7Aqe88XL1zRWK4Wqz8zjmPG8cC/cLV
jyhRDHFvZ01JapLqc/fc167Roar+Ecda6NJONDEm1RTe6KSRN5t+2iz8WqTH8G0JNKDSszIIkS48
mcoEnLpRR3s167g/GZQ/DxssQaiC1aOGsFfzo7cciz/cBMejCHwV2stJBuhVcsleDs2oz6K4skIa
OAGdxpVrXWvZiDqXOVLRe91GejdpWrmtcuzTOZsvhSL9ZZboZknMp9O2oOwLBpZdDT/2wU7rj4kh
vRXcyVuz/Jy3THp46Wg1tBgvfKjQcvgETl6L5HJu1iXWNp9bUtuFHR+opuDfZ//d++yxjbBn6v1D
zBrV7NanB3sfU06zr/09Nzg3/Oq4fJlnBpgTbLJ8s/wfe7wYbAbcz6MHa1AuLhCF0OQQN6aqpusF
xAD2Q/fCXqEUquxyuax76ZK0nzKLX5U5fcBhnP6bj1hZlF62coPxgOubAWJ6O6n9DgD6CIjiEp8i
V8ESbjugWH0iLa0cuYjifo8nY9WIy8+w8J07sVeCsew/Syf2NZ+qZxQoUDp7M6hZ++aAkU64WlCz
ZuBWrA3t+x0SN6W5WI7pMMziiVNiqqrSLkTsXMQac136gG8GQjgJn5/72BFfoah8+rLdJF9qUo8M
Q1hvRyMaLdEhXbhH/0OW2qeSa9yrgHyF0uFRxbqGPOlg/uOK8c4zSvrdg6EcQqAjDLm8r7mB6L8u
1Fsrs+1RKXn0CeGG2jFaYUsMIS+JGxmHYWUUpfF0HEu5KscSJXRQlxTbQSeiLgc0YclPMTIiKSoH
L8MSLLCw4aRA0IQuOwzU1I3yYqr7fcT3A72wbNXktPecqA5qIf2ABp9b8ski8OS9HfwRwsaa2HTN
EVDcv8N3V5Bq06i1nCPvsL0ckkWMCIWyPebqd3FYqmf7g0n7L/gAEDuA8xDchCnMXSQA5RRwaEqL
9YtqL9pfOOpa1ertAqZzZbeuBy6wdj9gjkcmqLm28rPXG6YioJtH0/5lOZWEecOVdnQvbw1TOj4q
vZ5igJsPvW2f63KO/FD3tFGS6cd0/cfD+jvRbLayZyiO2VPvOjRlUgFlS0bBuoV3sugK14Klv+v2
GTSTDBs6mNnQ2kyjzLvEPuznqZHFcL7aKq8m35MrPsU+efaKcX3aExoZuMaXBoV8EFgu9HkBybvI
Pg6/4uPZhQq9BKtlOz7B21ju7KPSRZtsRGWuirYDUI//xfeouhM+P2qyoW+6QqiOZEV8VuKuLfej
H3FUF1f7GaGucgF0ame07MdiaQwSJFxU+ub7nQ+XrtWr5nkQ7/042onJV1Dqbv8MCvbkrEaHiKDp
ojRGwixtNUfMxlAl23MiGZZ187UgFjM/2DKPdHJAR1+UXegyVcq1z2K/Rf4zwcWyrrvSgelAxRte
PCfs2ERosJqwQk0XV0Syo40f/Lo+7EPMXOdnFE6e9DoA/FFDYHPZUhV1w93aHFv0TjmjRbfcHwsZ
7txpd1s+GFZw8dBmYmgxJqDWFP8Cl0vh+zKCWvEUl+QB12GmVRTSNvV+l+3LnTxgCHGZJl78jEXD
Umk1z9AIdRcQelSfRhI2TZFpSzBW5M2a7ERsZmKrxsujdY0dcHeqzbSD3XAVAlDEPIwtqvtdc3Od
5hs8udswunBSOo+poEkbAKxEIm1BD1B5ISP5AFMaDEBaRMPvdmvnlovSoQFKmjXusiXXV5Af+HBV
1JzkAzTD2JQhNuXR8XQR33sBEGbZZOknO3B4Xyvv3p4jUAjaUEQxgFhpzGTDsEyIBZbHXnS/1frJ
/xYYbRAsSszQKwXB/PcdmSMSaC1L2pSkW63J6zv8X/ivycuFWR6RgvC3C/iOgT6BZw9K+aLxN/7+
MGSumjHQCVJpTwyZvl6cbE28Lg2LP5GopXD+nT8gvXARAbZCL++WIGjxzfWBMzvtCMi32xJzbSlL
N7W9IOGVYcOXEagjymNDWeMCyCcsTgQ2KN/TJgu2QFbUulqW4XDMipzbPtlZWOLT7D1QT8zQ/3PO
F1xjbKCexaXoGLVxSLm1SYpEuVz79oEizJzpvAIVKMpqzuBzr5KUH//xhazDfaQxmSVLOMT+nniK
eUuSrMW75nVu6nXmSJPTe6pG4TshBPCXXWzqhiJ1rxQAO52S/aSSf7pcfDixSVuN1EwaFPt+wRMr
V3M1AWlYFMlDWVsd3vk7DaUM3HcmG+X+1gL6Yc/c1ox33RgGIfOHIgM2xavPLMhkideGuSw7tNv2
rkti5+xcXTF/jmyA04+Y+0cmcDmRtHtW0LH/E7tDoNB+dwvT5e9HU4/dqJgkaSjrnW2ToGkj7bxC
Y56sWIpaZROgCQYrh5F6I1ycYGai21Cq+Qo6p768jKOhjzGI45LdZsHPoCZwcpn4ON3kwe2JUWhN
YupB73scI49JAAFomSZmiDsWT59q+50Wti+DrdwiKX+/kIikLyyqUAIysWhL3uHleFdzo5tVNnVB
rS+1ezRzH4Kqd74XcHVD7Irtdm6wveO7U2AbD6H9h0y7KAOlxxv7wPy6fkfjhcDbgEo0HwKUcbUN
2LHt0Hzk+9j5/gtOpFRYxXU5pYIlsovo1x8tXLkize7Q7zjuXhak76aLlgKj93MsKelq46XkE4Yl
OnaPPL+jD9LmirI0F+YKOSeQlB78za/juXm/zN6CFCfOqw2vabVn/LVGvamUH2WyJ22mSGylMgLl
LGGxBrXn25rMuYjO+SfsMtCvGnjXSnTg95uN1QVE6CD8SaBNRrY4Ri3+jE5pNh7hH7/4yKHxHxVS
vsBOH0Zc9FzM8Fd94BBAzn8Aw3S+9FWOomkqlvDyIOTHm2gn7xsnivBYhjIiVEPrLg5GdEyvWX+b
XHs8+n2uFdu3cbkh39gY/SxGah/19OZgIxV21NqhH+6mUz4gDUeVaRBZ4z6xD5wolpAsdh92PcQZ
sb4tLM6++wXo6xD0XCKCJjfUZq+xQkiV+vMkn7dhpYPUnS0J4oUAzPabNr7wWLn+h5kXR+1JkDwG
eH1KXD9c01KP8o8fPC+fkpWhJCYQCL3hfEImObetkixldYysgDf9pB6G6eceXPE9ICI/wCUC0Oq6
ja5ckXC4DaWk1x+ZtIf/+/jzAt1eIhim8lLmctll68NP9An36FxAHsHUPBX3/IY9ndH+40Q+pZIN
4ACfYe4ir1dZk1pIKz6NynByhhkwZHnsmwp/mKQ0A1DE/XxcXaovi6QZ0CUFxS2wEEcKWQ4e8bjG
SxGhcl8ZyULf7kfK/mRUwrATynjAM8libkbQtEQMR1w71mYiESe0mX2Mvp7TP12v494jaIH9qJ/x
MZvVpWFve0VQCdorLDZkmBMJGL1V8fTsYlExVieThwA9CUIA3a6FBR6JMVR9Iyv/GDkP3utnHqDB
js++ho7G1fO2O5RMUs8bgQnH9mVH3F8jwFnJOAytK2zK5DeYKIVgHmRR5C/9c1ZI4E9o0ToTAAgG
e90bBDim935D8+oAbmWxUCZfnWRWKjhnHMo/y4FfQIQC+SlfKDX41P4NcJdlQUiaHCaA5b7MfaeP
gkqYqpmmBagSR9mRrRWGBBVHS7NVM2bfxlA0HypiChYv77VXJReXuqFH45C1QmJGHwzNtNWPceZM
9jWWGKomsFQ+Qr/HAybAvEQ4dKxJ0RzYlyEiexhF5JGRvdR3tguOPYiPAGNJ7tRum/jZQE3JRgeS
Xqn5ZjEc2EW8fcLCL70KPhGyHdhqOI937uq8N3k2gCgKPDVAoChQ0MzljBNRPWFJKj5pFg9ld77G
K9UjFktlFcAjxlBXZSKe/fQxI44hbxIqbYnkVhUnJG0VQX3DCI/31CGo4/ZGCiTAh0WyJEFV0GK1
skXf8xX9lXCbjKowLgeiXQxopGSLWpuZlpoqNPU+LKiPw8rzlwomjgO5XCPIzx86ScwHLhS3qJS1
2psTkvAo7XtKqSolmmavLTmBgSsJMid63YnFilfqGUQ5LwswR/39J62iT08M8ATl3Tk/JjluX5hR
F+vQs3ke/k98oB80k7YGlbu3YxAYHokRsQZm58kRdQW57WpKQqRv3woLCSsk5oU7tiZPhUuublin
vCiDWfYSD+YEZFq9uyb/FWBC1eOKXSfdQVJ19QAr+JP3XeryLR9uXlbZWiKkbkxYZdBZkA7+p9uN
OgIs5rGWEz3eeMFHKqi5Jy+d59PZGy28OnE4657fgLXTG/7dYCtc2Gpk8ejNOUrJPqmumHHI5T1p
5k14s17oWd8+8dcWWKxgfcnZcj+gwg1GSY22lBLvPxrTvxkJtsBlPZzbYG41QO7NOp6RkVxUYXkL
xzlfdp05yO2ttPY84Yn8XkGwQ4jhLkkSes1Aor7kmRQJgQG64wwYHHQaaBkPg3uTNZjK0oWG9IOO
1e7Pjc/pRz3TTeBg/Xc98Av86C2POju5FlfdNR8bPrXFjXq0CSbZmcGnV5OHTjaEz+2QdN6KwxrY
2/iSERK+AHBiswjvyPv/lGqZJq6XDbzeUOibcliGJv8BJX/BzBCSx3OmKj0mJf6rkHGUTaRSgGtc
ZydxlUBJoyYqHDq9mFnw7EINyRlxOf3aAsB0+v/HXPWDTBpc0/VeAaTFjDhEOCad7LQJ9VLqQflu
HDBfuNtboCH18Qxs2DXl5yRk5yze/OQOkfOQpSQrHTpst/Ru+IV31n6ygekJJS8YTDha/V6gwizz
Y7g2KagE3luD6jhtU+6nzxbQiNxwuEo71wDALDSFw/MPjGHYts8oB7GvWbjJoJpk4Z+cUfu9J2dw
ZlkuNMDYMayMd3KeF7xljNuu/IHHnL3DdFIFzambBm4S8ivaLturCiQ0w3kYTIJXnM4aWfezeNS/
w8WB7vGmfykNUdoJBdESgAi7FuFyLWrvQb/S1xAgGNHdiq4eETKg4kCES93ZcBS2hv/gpMfpA6Rz
YSE2xr8Q5kO42vThNOdsBEcB5IP5TP6hLcyEOpQpRph/bRpy7hZ1T106kVtceCxe//toUIFSgXx6
sQmSzOonSj6fDj/75S2HXQju0dwgk85Y0nHiZc+f/iIkGfC4cageVFSj9CBiciWInkdyO4Ne72AH
oVplvrEJ3m0vCo5eL5veWUoqnz1ow8/o7yn7DRKlnHJ/oluc2FCM0yT71TRBmySItKVLaw6IRCFg
mbkkmsxjcgaKBtAdaWDw1MgQADPQFGORMwAMMINNc6KmWlSi1gv9n14Y2q+C+uKAzMAmi+bURxpZ
7rm14ic5d/XFDZbl3ctqz7mOID7y78fyQKK1LrJbzmJVAbAqL4u8zHhWTP6tNsoqcnFhVblVjyKb
Ca77tTYcp0sm4KvL109By/MkjquTv/ga0QKRFds+YAav+leFVUwQrIFdxLg/s1Gw7261Jvo0qsVw
Z2BbxiNkPB6m9QxEOPA37EAS2otdalZIeWuVmWa7S4FioroPuzxJ7yryC7bcPy6mNiiZhaaG4o/y
tKgn/OsoH4up7Wfn2dhGTESDos776Xmwd1xNpTzwjfRAtKLvag03waRjihYnD6uLNuYcb9mVSnrV
WnMSoPKcNPkludqQCA7XiMeUS43LxzNeqkME3Vdtu1klzsogRcdZLPtmLWx1Q4TSS0SZBGwmRwUQ
eecS51TpDYEXIvvxOkhz8w2WxC1z4genv19MfBqFyOYuySEonxoCkpxBUpkBqcpaE1zDseit02GQ
1gdJ1Iyr7uowWCnkX4ddfGyZEqoER3rmSAkgepsMJ+4p5lgEOdMbM22knnMdVY76rQExy87qSDr4
vQdzMn85jv4NWj0A0fhZOwUDWW00YrOQnavnTiKKGrbwH03mCDPxmwmJTO4B+9dt0GDMnHzSsptl
83atu3Ywk22uZH0scSjANnanp+P57MM0K4EtB+wFS8vm6pYl05DACh3WPi6n++LTUHP2nT03OQG6
Zq0fU1UwPuNLt140rYoWyXo/R66yY94g7fHu1RCIiKDkder4mfpRpOYi2C4ERw+wB/uxFdaFRxuc
xqx9cE/YIqs0VndsW4MkAmnNzFLxAL0AOoQZuRatjXwpdfYqOR2zAknhQPnDfv5ncRxk3b+VFfy5
Ow5r6+SoqGEtWyvtGk9vFHjWnoyE6ZnPHCyzH9Wb/8TNjKLki1E9Zkm8r6/HaPUMlnVrDzlZXTA+
l/W76ByRgiaxwRwmFuhqsb+3eO7lEGTkzoTzV2Vnq3mXTfqoMhwRrbs21dahe8H7G7Q2NRUAhfjc
8r6kdwSLvALjsHb8+7OUh90vUXJpmYM5mRMrrdODavhMDoCmcygfdzao6ta3zoYSsPCClWWvPybV
GcBAJsEFTocf9rk4y8UEsQUU8BS8xia5t+ulPgYQx1TRvJNMVCU8c36oEdXDuCEL5Y4X7xkMuNyk
ATCXGWcNo7V9P3bR63707+nzFduU4UhFf0h5X8AcINLGwBx0v1XeSMKk0Ym46oiOgVMeHwr84sWW
dd44Qiukj9MSWMfobV9FiNBLV9CAAqDKBX3X5IY5M5o1PhyKlRxi6CoQpvqHA7e5xXODMFnKvsbD
+LQ8aJaiOp5IqiQYz3f2bWt2k/WyD7sLE8Zo7mTwbASknZjSjkE3xVeNqd6NTfK2+gcnUcK+izou
jdlWqu95ulojQJxFmShn46iqxhdbxvN24CrxOIGoT3yfkk8XxfSbR7LND5XSr25x7+hxF+6s7shj
j0lXe+NQAkGpmPdFVo64nHkhbdzysHQ+bNs/lT5fuSGrcaFWUB54JjgX+KhiX/4hn++yZFfZqLv1
QARi4ygLQSTmmItDP4MH3LbZK3vK41HJIjExAz9BpYl/Hj3+2dsRzHE/mrou5K5Rh5efV7dg6xOr
FkkWfaESOeSK/QjOv3QUZd9b6lxELAtDddYEQA/0tyoWtC28buhcoDlm7VhwMckusGQ4owYnEpl8
GMd4KOoA8JY7ovO4hulRitb1mq+C+2DEOZUmni+W4DjvhmEGH0VHzVYRANdPoT/5qsd38OLZ1Hj0
E1v7RsPXgwEr4I/CQNWapAftAshRQ2wo+S+ycFmybqqMHz8vQbpjdeMRMtCmmUZ5i5tp3wLR1U8S
ABLxRdEAzLC3YtkDgScSli30rs47G5CaqjsM592DhE4cFQxAwaRawez/XivvwesRLzdj873D/Lwa
9oqlQeBoG+cH49w3acEqRwHLyE7bZOmSedXAFdP3ts/aM5vEpOhTVmyGqLRWUXhaR2bx2DrRihLF
LwX318tO71MMJ30T3lXJKTVHGDX1QdkfMLua8wFOCL02JW3jMaeKsQqmX9f5zZJhRWmw7+XdjNZp
lfbkbt95X9Suiak86RIdcLVAkiI4cwK2WparVpcbFck/PTMGdMOaZztzGWEt/um7Pt3XN4Cu35Bo
HC/4Yfc/q1zdqgtblJKtjpnIvMfY3ICti/Cl4a+am0VkBXJ/h7aPdpK/pIZK50F/ZApek4Gn4rJF
4DcqVVQAfBMm7sV/WU2UTWxyh6TqtZWZp/T0rS1f8f9ILBGyMGbTKyHFhyB0Gr5dNxZNKMKU9Uy4
8AiKxnQxtRZFpR0JFNEufp6l5kMjshTwFIBftA07DxDS6vv25herpIljN+XBUH0c6cDL6KH8sBWD
DAd4/2jrrXpi8C/4GKPL0Yib2FgyQkIRrI15SUUzoalw9BiVF1PJlKoEZhvj7+rvuAQN8jFw4ROF
/+Q0wI8CUEayr2srn+AQwVn+chlRI8U8Zz755QwcDRJM3KmJbKSY8cxaFDdY4Tm+FKaZTe/Ww64K
BV6kT9xzQkbqD1DcWyPDz27DpzuyDBpn079oiIfBfZFmNGScPPrRjviQY4zKz9uFQyN0sVPNKs7f
CAcV13C5D7rOl8n1fsZa/a2fkfZAF1Buhk+74TOGtZWSXsPRb7Ud6F24IiITD48SE0jtq1H8BVST
WEzK8PPQb/C5rBPPdH3mKj53xzFPHa84Kg/9hdbaVWHN09MgzVu1KgjgG7ZBlTJgu+XS/3hAsFiX
JjiHG2EmM8wuyA/XAz5G0FY/1brFofEn5igZuHm6kpE/jr3KIbOO1lzCPIzS3gbRCLMWqrTEXhhj
Fl4HN9Np49GtZZK2CFIBmgG5Sl8sePZt8WLNG77UO4VhiSI/ZFZRr4AT9UrWSTiaPuUN0qFYFv7z
Ib0qoQghlKQkpDFKGQiuWgk61m2Oy55ZIakwZhYjPixbeSukEbooW/uAzSURjjBJcJDj2kbOhFwT
kcJuRWCjl0tWb7fPGIBECWFA5GxSRy4CV6pBY9X+y1nwk2JBv80aNFj0H8S5zpMEcMcD9wzXlnOU
OraINYhNMlI7pxlBd3QT59+yncSaoIfB4POpwy4/D8dDmIkM3GvrhkwDlrT8pwrNm/GhtClcAhAT
ux9m6ZuSpBIl4OhB17iJ9qdgiex3Bvif2BeaAXApdlgLhEG09vD/IMYfY+QIuwAcNDf+ueBobcEw
LNgID8dMaYzm04qfQXLhIKzv6wfshSs094SzhlJew/epnB+NsrmU/A0T8dK9R3JAJU7PPxXWoG5N
cHaMKf0JBkFZ2v8wCpHajaaZe3z/MuLv/WmcCeGgwJtv5fegBL4hwDnfywceqWbiR+BX+Gu+lHth
MvT2xgc88THQSeQnSpzT9oRpn7yU/wVCW8Sf9b9nJPNqNZJhwuQw+JEtGR90GItB/rF1CmRnVipV
CVtPQr56spDztolMsvvP+2vK9VjqELsYLegDPiqzgIq+CGaaWWjJHjiRRe9TX6OHaCZIs1mELESg
9t9vUGKZvxdOM/gCm9ul4gePeQZD0Epiz7IMuTQMyHmW8mhf339Wg4gj+WNl6qxrdvOYnSoZEhN/
OWWE0svjh5t37bMRScMYUik1p0lMqLIqMibqTQmcnIA2LyK/jFyX2L6ZiXu49B5osVDrUfiKY4uL
bgmHtkpgQNnuV3Ez8EyTCXdLuce4Pt1JzsTJ/ucmk9nwPeoZurswj5F06YO+DG/i+7P2qOUyqsMS
6/HdDvwP+Q/m4p9lbvkbF7EKBU7vfxJ7LiPraN51UGXZbBInhIQHATTfjqTu7TeAMkzLnIY/uyf1
axBUr77P5vhaAObAsDC2+x+Lt1336J19ueCZD/z+42A3cfNjkqhgkVb1+XT4TyWfeIpsWDdX9YIT
q+gMot7wUr167fmLl7v/6S0R1+xdNgJdgr6Kef1P+Rpvt3ZzKkRVsY38pXvFrff1r2kNDiu4VWU2
M2hRRy4zRa595dT3oxJhrsXiWnd4OBb3WEBvb+CGTA0S1VgPG8aEeYri5MRKP8UdLKtddbc6LvnM
bONhALVwrHr/NllBy19vJjojEmVD9682JHU4tiQgx0vNbwl+mSiQQS0P1wxJBeP/w7xALFtDt5ue
eQO5y0BnCMT4bxCr8xcwzc7XXWegIID2uenEd+rc0oPSRa6ZwpBAQwtiBcsEjifLzylzwnihQscz
A8/WCSYSTwAunPsKwrptAAgaI8f09F/WbyJtxD8OevaHQtyx9VZW/NOX4XtS8EmdUCKafosfiE9t
pTnRxsMxYx5Z9Np8pi2St7zMk5v3YCBgmd/CMlxxBOwFOj+3nv154BxkWEArRaaYV60c42m03RkJ
A2KoeOFjFaiWvi+XO9q3IWehITyxTFCWSbJHwpc4LHY7I7CoBvuvvqCQbHm7v2IZGRf6ARArujZ7
Q5MF3fIO/apV/KfwO4GTYDMuQgV6ZY5uicUhgIxpPLt5eZZ3zP7EaB6phLHNp28YR09rqBa6qdHH
V6cZeECuX/Z4xHpVuBjSXP68Nzyjy8XwTBim8sJnSU/NAksg7FVVP37kFBkf+bIfccnHggZ2KBCI
OVz6YjGtGsJsCIZWAETiE51aIncEq+BQEm85hL+PTZM6mYjmnuYKDoqZPWoHTE22lobtT5KL/YcE
p0VK/BLTIR/dYEsVOh4Hq/PUQh8GYDFv5bvIDLa51cOe4xr1eVMwqca85iNINCAPaao0BYABQvvB
njyMS03OfMObvJcKTXoKFJOw+ouQaOq78DQiljLPtE8sUuQvWJJV35yek1rDCoDXwcnGq76ZCtTg
xXfjxh4Wl6iDWv+FSPRssAVs+Z14LHmuteJKkAu4johJMmWeEYkVCL70whsIwx9pQteyMpVbIXRa
62rpkI5Z+dNdvSPx+MOy3RFRofLZQDbV+Vt6zbfr1qi0yqtkmtwTT9Fypbtxwp3o9e0IPelO6IPN
xr+a68JqK3jiPxK4knw4w4Sp0Myn+U46XJVsoMC4c51OEyU4viiXswt6nk9bETq3yAd8QmQSwZcN
ndx4+ORL+L8Gl2lZc+r8CVexmMH7oVF9IXOA1zM0/x1jnUUl/0Epz1d29ECfSPVOeEUB3j3c1Cvn
9bs6YDUef0HU6zQ8HgyMijTWCJI1fATH9ueZxAmGr2AssWA4374wWu+qh4eBZHjD3T0TJnvDA1EN
AMNQvxg0sEM1WH0YHbhjcdapOXPfk0a5cPzVVJ+Yrkmf+AOPUAbRHlDZqGAIIrpx5yAHPqJUAUaA
StJwItb4+9CCHD9MbHw9dkJrb9o4R4A0wMgEbtWmXDtEZ2UneGzxrgKA/p6KB/bCm1jiitifdQUo
OYva1f/Pg+tbTAmYTFuMZPgOGERLEcd620WRj3fAbbNvXLASNSYQjVQG9RKFpO//9+oPtUMK9qvN
RPETrgEby7U5X8UvY7JwXhyvq3FejgxFh0g7oSJiO3B/BjR92nXk/tFN7i8bydeVn5d0H55mZBQq
uVyDu6JtVscnbUXG4iNqCcI7xjVDkBvTLYFgLloeUFOdUmKTryO8+MYjGFGph7Vg0peM65H3toqj
fEZQJyjS5GbYiAsQSCOpU/m1vFFEG3hvQcnUlbFREZBYEPCm0do+9zqwFPekTyq18Dr58ncvFMSz
39PiHWc+0n5Nr4bDWenrU3jfovMITfqFbwVXVAPIdnQfRtCh0HWwlsZzDgac8oddmyRgo3tX9v/U
QhnQ2ruhMwWYjLX0rRj9eOVw96h6KRVdRJAemYuo3QxksEttkoatZkDHUe6xMFXFgIl81uDzO12w
+zV8AuS5MojxtoyFHnc5FTvpVM2dNA/uOyQgYV5GqF0OGXlabuOKhPNlbgUYTf6cWfdZ85+cv2XT
JNtsJ4H7/2/9tHW+6GDFnNkfrpvqk07pnky+G3xXDjV5SLMTpitP2Qa75GWow4jkxozZzjkPiVyE
TcEoo48OJ1Np9a3l7U7DTcRnbuy4Je/aBCBaUEoRwa0JDMrn4cBPJ/tpbshkz+KEGn4+9OznC27K
3wUX6scxW9iKsMEggilC2LNwVtrU39jygc9BP+dgolNM2FcMWP4k+R8xMBN8NPTsbzIgPR0EyjDj
wUef4sqUJQhSHN+9FuS6T9t411D1lQVB+zTpeik5EscDIH/7F/2t2ilL8CyyPqC8Wl3Nf4/PhjAm
PQRzWEPxm+/+Wdp6Q8lY2/56yML/9CI+JY8dv6SzktjaQywGhg4UbA9OkcE40v6JWu7KNvwCtV6Z
ih9qVFjMUgdgavflpQXK90WwZlLUuQ+mrAS1CBsHvvsegPdbS4r6QSniIdUTWlzdQDHwAULjpPNB
HLOaGaWgIiVPIo0XAGDVG8pZYTruBnUgxgzWEPrWAeHXiE55hw7bothB0B1fD2LIsAXW3Sy2J4sE
P2qIVybtsytT+i38CDU8/PLQVpa+cDCiiONM/Xesi+reM9GM1Qn1dZuQz03ovOzod4crmzivCOBO
tgsUGDA6hmJHxrtlTUJlFxg+hqL/FO+ZkgLaonidqfqEHoqYSdcNRj0Uo1ZwRZDn9N8YPR88o7KF
ypvkGU28Efh+pZeEpUgg3k6yNNuO3lVm9TpkCiwiaRg6msV8xlteGu+DzPX+dreFfbxSRX0xtZLi
THD8jHB6503LlM6E8CWI9S+/7MhgtFA9je09f2TgkigEktBk/ZSHbyrZofu4pO4Gv/sa7cb1DSQ/
mIR++5VobSiRSjD7mAqjS+dMIC548xbMqcvGxamSAW61VW2J0nwVR35cFW6F0/aMnH3b6oQkJ+8Z
LViuWJbeOsz54o0FeB9N7B4D2Qn0i+KZNfBPvfMXPTrf9TI5nUpFUrDOeawX4b6GDvVyxV9U2FPK
ppAnL7cV1K857DcGa2jFEK63vlNoj0AQ8sxRfJc2zXgMdk4MhVj11qCzpaFdidDllzFao8OXZLxf
EN7Y1n2kXfJ6Y05qCMd3S6FCqWjYvXuGTjjGaQXx6Ghb2yWwqXn3fx9o9yf+6I62+TYZ5iqfX6Lo
UvTsX0LDn329lP/znXy2l2H1YmXI0nYjqsdlm/prdCRXWE9VqPYJ6B4St1HMPGzguNrDST/2Dluw
1n4luuTJGa7TDbnzMGK/5RLheScXcejtJAdAwlygfzHx674TUUKbh/uEur9DmA9H08e1YCojfd92
jdjT6WyKlBE2i1b2lmlTRVER4R2FvNK7sFZVnwAFLtWDQWge5HZpEDm1K5kvoWpcpmep2PayWzYo
PPiSdwtQcRLRE2n01sspFncx4tCLC6SJFvGpsDc8D5zIRaLg05xe1LiaBDanTpcpi5YdqH/FyQed
bPhDTFOl9buDVNtUC5pv+cXy3rNtJhmPOmZUAzAqwLysBm4WZPSYbdvktr9rKFEJ0xuGAJmbKzzE
mtzTuLBwxubCiJWlE0gR5vsEXMq7Q1fRX465LFrkHhKbnx17hMZD0BsntAzWzeyooAh2saNu2BqJ
z6UqNGMdbVJq0eQx5W/+BNeN1d6OvK12F+Db4mf4R6tsIu+3gXC9ILI4qwwsYdbbtIFQb7KHd5Hp
yrK9m8eilXKrMLAoMsrmZK5F+juZPYU7Sj2o23/5ks/ZZmZdBZ7acY2giYcG8uIrTfxj+UXQK73u
L9Xxa9bTTgtfkEiXuFj74SPzA8bB61V8XBrQdN0RNxPjdpEtSlwlkun/FTpBMX7ObnfusRBULFSF
glhvfxbyTxhyuNwZ4L00e7kPWbY+jAZNJHMY/7k393ZxVNCfJLsKWZOiyMQJkCJIFqjQBLvrktc8
lhUkueqNLC8nnED6m8NMZHRT4K34BS+9SF4CwRcUxCh0FqSyIWHvX5WKRzvo9XzMz537/K+dA9H5
xLDpZ04loXU2R52DmuN0laGTXwS1AVw4je1QzRmT/+5AiRiKZ+qfEldFSYfgGZqLs/rt7gz13T9+
B8inSgSfvB9W65Lrpxa/W+gSJagTMAZdHCt/U6jN3jPP09hMeCX6+Rr9iSz/5Curq6SP662G1SfN
7KfTzFohvwuvU/v2KjEpIeeygSErH3/f9K4foTmglSXbbpYN1T7LQRt3C6L6zGgaeop0fub/PALU
5u25P6OHobOLD9bVsl1J/A/oITNhn0rZamoFGgwzi/A591NNfrnkKijKq/PfRmrzr7G6xNVQ5yOC
sI/S7sgvWZFNpmPTnzzCQ+affXsOLroMvKeEL2Uaixqj3GHho5fi+af5aGpTw8ZthfOUxVrLHEpa
OmFWKoGF8p5T2a9/7CJinT91X+/vOjBSNbHROqLvOq9CZU/PSSWnsUZn0SvwdA4l1Q1DkfdZHX9G
jjzrNLc9kByZ6TpEAg/HWlaCLKVzOIa/YJzEw994omRAXmE3YG4fZtOv+kv11eD4K9JKZmMtQ5AD
3j/aHkAuDbOXisTlcmihr79XdVfDppmyh4lqVw25vpIWCGxfRCN5bmu7CiywbhIQVcP18vsKsQYM
vaCV4zEI2eWvEXejPfK5TGcri1cob7OZVx/lhU9vvfsv7kA/VsFge8Y1Upg0ccN8g9AVDEPh4lKN
j/CegL8CzFrG+KdR3SJhEAYXBNg7nee28ac4nTAc31fHDEJvSJYdkb2EYNh6j2pFF344oWbSQ3m3
b12MtkC+j0uEB0CNdf3qWx5epqhFfyBRe4u/GLWPKRgMC6UElTf+ew6zI80GuRwOhOK5TYe2UUaW
skSgq98svhf2HgXvZ9SsqUZu/9LfC7BHqAUQsSb4nSpy5g8mYRwwD7EKPFcC6xR2oR63s7Z3xp2O
dMK6JYcipGxNS7kdXTw+DT/IimAYr+AYmJCWeXqi2qxUnYgLBcBfseHxEGYkeoh8oZXzwA3QF3tJ
kY9/tQiO2KT3L06kAahd+9zpORPhT83FonWm0Me1rdGZcUSmTmVzLtGggZMv2I3D/Nzo441RDwQm
UqAlX3QEJAClciKFEtXcexCGHCbaPqsZa4iJ+fU+ewJtMxsi7cFHRQNe/H+Qur0G2v20p2mGd2Id
G9AWLEkJV/xp1YlduVttmqig2f+TevIETOAqwUKAIqOmy9Ws5+hImhMOk7/ST29aX6A4Ocw22o6m
aad7Mss1q8Iof1hwB8d6Gyk9ZlhniHscayIysIe2wtTiv8XWWcp+n1Gu1obiTH/DZr6/QBrEJ2RV
NNPQoHjztQJPfzRd/5FVuONkQ5WIGjXTJoVAj4BpEks9Dk1E1bDWg1FunbzbAywmAjsD06R20W3S
BeJtQLP2EVWHyhaTBAf2xrTI454b4S+9wVrUJPKiun5MpQ0OZvqSIggNZnGnYmB8PK5R1Yzt0rj3
EuZYL39RLCM/HQ/KzwWUdmVdBH2kFdiyK+OhJNXkYhkOzl8CHw6/EFj08WLR5hZ4LyjctJ5x0ZwE
PLhwkLHJKL6+YDwCQHfE41KdXLiyzveJOEa22AH1yO4ekD3Rn7D0B4QRapzZ2FopHXepEWvV/Tjs
jfzYezYyYcpHH6mREPD+oq44GoGkRKKxYOHamKgR0mcZT5218kyVbfMAVovazVdYfd3tiJbbURKi
9ZiA/Ycxp6XJTD5TvuhKnht05MCJB3fqaQrVsFcQeSYQgEEgiHcbYRpQhJbMKiiphlavOwriiuvI
GxWz4YBKvEaqINh1w9GWw75podPrgPIEVIUzElpcU+t9n2OhuJnDMafvTPTDc1UuLVZKFpCOXcPF
U1LCaxlrwQfkgJ7hLzPFzv3YMfOJtMR2aLTjGU3y+LBzA5Z9LSlQNqMaISj+/1Az9zx8tdWEiIjp
6tIOGxAjy7Bhfsc89zyYrteITFYWWPw54DRK+ToFqxIZ2fkG670qX6HCQCi5bTKSMUWYYDvf631n
kD1S9sIA2Nf/ccxhP390C8gxhLkKZuzmPCpVwQOvuqBkVoo+FH//VTf3dJTmGYiE/YAXts+Ih62x
Lcy0151Bv7L6uXxWqWzP3BrEvqpaMXsVwfVGxw1W0s/xKL0hrV4WtuPe19KthGRvNlg/mXrvM/dM
5pVC/2PRY8rbXswldCHkrbHtkxmbehMtziK966LxzpXFIJoBewm4QEJjb9M0sLudWyuAPstKaFrH
oDI8DGy3ACLnHPApVLw1iINo7Ts9EBmVc2poqUliYqFlNCWDiDypk92WE4MOUz1tjU7j2MAMSuz7
g0cimZTZ/PB5iSniZUejk8NFTa3vq1wQvfsqIoEyC51w19hfbKMsOA0PIYWq/X/LTfPK/cFDW3ur
MjRvH0vwX25lIywZcZZAYGoxQoYfq/8EcMeGHbS+xS+jSLxq3iKvlzba46ZvV94Cf0seG++e/r6t
Y4/4RJS365f05zzYwq37ZrFW3/qzr3B4ci8RwJJfuAtd3JGE4o/bDPfOYkWtMK8MILJG80sPfgvZ
hwiVixq9MdmpALyxNJKX4oZGDnbN05Qa4DBSiGPPYhXoGRShrTL18hbN8EjJGWLM/zSZx1D1QpaH
vFk2+Cp04aD3iU550uUQYs+6uLk204V+YPNFQqiH5DhWUA78GS3X/66Zf5tYfZ+HdbucI+rdF5Mh
PSproBxRu5lV0RqmM1Z3veskMnsiGiIZEvkkVp8dNHtI5T01CnWIXIWHg08ySIHu2XDl+ddwVef5
SLNI5dzSUn2+LHMFAwPgcRq+LdAL5J3kI1f6I88ld4Jr240GUTcQy8NKsRY5oxReCLdNWVAMDVem
nPzX+4yZhWgpFrZ3YcDx/PZbXxVNJ2AoTjm0UPOh1oADb8sqjFCivQqIlGM5XD6ZQ9Qgq07ftqPk
/o5XlJFN0mrZuEYbDZbAl2Bf8sPhsVIcKx8w90WNmAP29f6tIA/QXtLUO2eB43UBpFcB2olOTO+F
l+BJxtBUkvaJf+ow7A5ltHReAvQ1jR8cGM7dgovLzJKN12NgKyl9p6s/F5chDm3Vow9RkG3TQAZx
fCjnHKvUyyzuUpQrwoheLgvmYzLOtTYDCue0bnwQFZJHEYFGIFMz1ki4rqAzZmFCVo0Lm7kjiBom
mDnVgh85dCNF5GpTaHiPgZgs6EZ1MOGh14cbWia+fh1Iqtoe5RrBmJ73dsKX6UOCkgVlvVZ4zQQr
gOhMm43HVyMEZpcOZeQnRudJ619tK8xlXAvv7wDoQv/hA44YGkghcIOLqRI5dSWME2vl656BSE7e
5gskN9qFkOfL/3ncYwSdjRfsbja17OsbLedgm9B4l/Ru1YbRdg0nSOEZhq930dSHgzXTe67fxVno
ziIIWA6XhghElf2+r9/TcNNSMyjocSilrv08xWNZzkWk3C8ZkYlovbFhfqmTQO9xOLD0kEqobNcM
iujS+8bVHcQmuLphHYnDwi2mtIxxLdBsRO8mOxp6GpPBBqYsZft4Bs8qHsKtqEV3N7AXoeTni0qs
/tKCUGbm2JfS4V+LzU3Uq1IWIu1sJ2kfNT767wtyrmSzM0esgptsFAKftblReSoIf3aESgi8Ns/K
7Bn0tpsCvxymnD0QmgA8xjByYiVYPbSLgIHQKjcn2Gn2hB9kzslYawGAWUpw3d9kdubAukpr4NRE
gff5y+m7LdfZegjeeFAVVY0StqrNcEE49t21r0QKFVFkI/p72QIxqKb6zcIRZDviGRFWMvffh8Go
LgH1VYFkEfK2ceAj0CPygBc8LzJ8USENQHCJS8Wzz3oJsc2WHhJnrwW7ZaTzwbpsxO/A4xHTE5MD
CVHECz9bv2Ryi3LcXoQjfRkG6MJbNzzusPXqCusV+slWmNNVov81G6SkVylE/V9M3LdCtJdpU9dP
h68foQRqb6xf5Ft/Tx68mMPIdgbKxZyQRiV8jUEOsMB2zhZEphbLo7ZvONOUbhoZ9gGULytc/wEi
QYUGfhGGtxBqKhxYdth2HBCD2MC3SS7XsBduQ2aptxmnma/d/N3xFbHLdfX83zqQiSCrdwKAkm5E
MKLUegnMS6DNCPiCqrlxXDxg6haDxDEozgEw3fVX6z2/VLB0BuRMzdaxNK4Dnbh5+mn1RD21vjZJ
kix6IJvzvYvqhYxnIAVSrZ+I0yfw4DQuLC9CUQrQgbFs+9x9/ZUF7VX3yBUoNIO/1raHtAgnkKpC
0aoHGYPLRTvnCT5dX2PQ4CCmZRs/fLJyRKITmjLN4yAybC3r17XGiC5pkT9JavwXcBolS0ZXitkf
JsXr/jHIfjOllJVGXmnLPQ0bUt8ReMWOVQC/V7samCOri8qvkjUQw167h3fKNT7r4Jy8ZpRRV5Wp
Ffi8wlq+iXRzyTGNJj/c/s5W3lk/ePmDiB27fqf16tCb5ie9aLjlq7zwAcbSohftgJEKv72akFWD
onYKfADfOlYwoxwDnz1bZznsd7bq55tF0mfnw3ncIgN40q4XP4z+2jIl9tcNIv7nyKtZ984Ldkk0
PVj7NPqURq2O36uy9uDglZtOsNsXmC2KhIyJgV2d+9XPLCqCDMRytalv9lo93+FgnavpO7PXBBdS
3o3fsKZLjPfwWvMWMbv2GlPi1rgXNHVutk/wZALj7c0rzttd7kgRwcbhagh7F2f2XUzSnulGBdVG
1gkqYfQ8OcXDh9T7ZRrnE/J7pAC+PFegvOyFP1dL5fMy9AnEIHle5bggiVWeFDu9h/4KkkOzl+Dm
AFTr0l95l2+SM5tdN2Wx+DEjuynYhSGp3xpQOuR8uUdfUzg0QoEX51YKevUfbIVe77DD/99QnPvm
jBpV64yKC1aMKpPwc5CYIXHsP9FDzzdpqkMSVbHvXNpa1kFrAjg7AHdavc6mFUknYLxS3r7baZdQ
KNSzkM7D0exHkuhboMEt8DPO8uYfEGkDf3TKVR0o8sNqWphxwO0Oo804ZCudCbbq8rkw1xikbUWY
w7mAUsNC9APCn3ncNSWwE8G367OfMcAdF7c7x3cADZaAKMEM4p/aADWb7oWdQTF0YlFdm5zxBPXo
klL7gdGbcDs+1s0MliRMqa+czUY34Im0YmWAb9h/nLqGHfwp0Wnzkzd0IfeF8eUDzVIkEobQS5ET
bNsf+3KwAZ2j78RbydNwLu+/+/PhswT4K49mAYL0/SDw1W1nNBGDXlJXcTk6svT9tQvfDZDmNDZV
9jiywxCFyxQQZs89k4Y9CwZyXWMhAnI1m/ik4SwEIYoBwZlkz4KbR7+MZMMKo8kuyD4rdDUM2rx9
rruLAa0ZGPXsHGiQARreENItOtTPsumBqseCW6JivG8Wzll8NsX73BlR11ZMeqKqBL17jL17Kaod
RHUIQ/TriVc58/np47MMvskgWx/yu+8sMjkfgLtb+GHEmVetmhD4fKMI1LLdmuE5DYDDOvXL51cu
wySqZ4a6n2mX+Vt7dxW/VCXN4XPHLF2v6vYpP2DnaTWV0L8LjEvpMcj2n6K/+St0KCznTEKWNXtg
lV2v4GNqoY2h5qtOxt3jIMH0VYPcF4dKZtmssJk4Qna46G2WNKwQMZ7Bu0dg95rlmWrGcK3GKneU
y+bRmEmPJOZs3KeZ6RDlSLr4N83GAz290jRyxbDsMK5GtPLZojvfxd0bRdXv44Sapa+ULECuvfmx
wtRWe8DmBiJqegTPyWEVK69rvQmg9xRp/7RLZAekRv9b8dJhXAtFGerw8sOUW12oYKQS+vt9if9O
ZTgXdPTXQuQNGZew4eeapDMltaUbBY2Pe6Ykk2ACe6W94mI3O/ky7zAyJkYBb7MVZojjIT0r8Nk+
icJhxyi1LA/jHqfHxx3rHtrajZf/ImcFz2oiXjv1gKJrSS0VzsTpDR3MuOJT6dB3vHltmNa6piLo
riux5IvNTrovPyKVrlyXYFULTkmmyToZIaKKcxzObIpSYILHdBO7JL1iqAXXVWwtJz8cXIDa+mzb
Kc3Cn0TlKbsg4ZvznBDQtdYS57sTKPmI0PioZ5EJsmnbThJG1wPJGabJp1g5qPhr3/RKbqytP6ab
U0Lzlqyv3KN9wT3IXQEmKOnedNdSWcLCSEa+uA6ogHnEx9yyWgwSwX0ulPTiTSg4wdaAqzCqYBZ4
ABCA8aHbUyItggWmWwxE+FS7DwnR7RlrCRVNrGu8GvTcVpySnlpq/GGSJSqH0HPxSbcIN/kP7MjC
cmC1aDPFXOuHEl0iE0rufJO932bd5Rivgb2lBY8VUXQMI68W2MHl6Ayaztxi3okK8XDGseLfeh/S
BqutpGPHIw//drqZMUmRM4aLtLxbBFlpWP5EyQfu5zERdJ02nX9M4X2E/pb5VRSbXQI+C3RNvFqR
55IpRQq4bqkGXX/qDnmOX56QmwyrxU6YmHRsJJiP9xeJp9PeXTe/1/NldqnwRWeQRH1g7l3wuLh1
99O+Prw8fsTOx9Cmvl3j9QT1/6W+TvksI2EKBSRC8tBVcnaHbktIprK/+1kcXYy0R+radBnK0be9
cqZON6rfsDXE5l8wbdFBHd/K1MTTalc9ho6/8H6aMlkB2/+2mK72L3gLZ0zd338yTASsuFr10yjd
RirCQRFFtZCvxOMuH6wOWu7U2qjGB4WriaY17wdSGZYJsVGcsw/u018+IV8g3e5/D+HzHzz5VbAn
LgNIp3ecIOZa/g2ls0a/AlWTWAKIjfJmPFfZNtSsOA7ZGsMzZoNhx7GDUHNafTJTgw2VlV6CFKg/
L4BMYtq7NosHZer4bkdA55ySdWW0mY7ycI1eXEKmbJ8EsacmMZZa2NKESOWXYRIsPN7VGK4b/g/6
xnohDO+/8O7mz5TjRAHukpxvl6omzp03ZOvJh2O4KX7qYSPpmQIMk6sk/tCwYtVsi41DSpaOeMWn
4A2vKtaZ5if1PeCDu/fWCvz1XkUC3K51WISLBxTplKlZy8aVEWvEaPiAYj1uzuYWuHOuGWfUlJWq
gAp8+vT9INt2kM65FNWBfSQoRWH/VlOmHBs1pE/5jn4t4Wgend+1Q3qE7knXgPvaegu5XEtEe98n
WYcYLRu7SAQvYFz2VpW4S9SGQeeYBVonhHKgEzjcADt7PO5S1ty4KbkfSebGjINlyPQQHpDH8Bio
MGAPOWu6MtH51bJlzMwLipvyMCzH+q9syCVYM2amehKJGx4YQBaH9Qp/lhYq4qTiJThf06Jlwhjm
HOkWh4aMg4xLHZR/fa3RUHbTtRFW/Uzu+gMu+p8sZCeu2OHuww/2n9P6QxW/Ny+sOVn+uB2dtSp5
T4454559qX0fA/GwjykCcITba4zbRbN+NDytncm/3q5WBVKWg61t+itOhXiisckyN5Elwk5xuwhv
zha6uULJsQBJT1zUqnuoonccELAP0oJqq5ffkRoLpgJ0nm+ScdaN0q6HYJVCu1Eztzpt7KH5/Rff
yitbpPJWKxrsoVxO0F2rIChTDHqJuqpFVLkv0xMZS5UhF9uzi+W/541Onfn+/kWtsGGE7Oyr5iqc
PdR/CUJKdVB2c4w3KEG/onExSeQtVTshXU33EFC89oLIdhvb44X+eSwHTefmB2UKa4NymtXCKG4R
LRTKegud6+oGRRBE6jLeDZbXtVOLndNUzgzf4n5w/2V70f+rvk9+o30qQp+4OhY2NHqqgVppBQUf
ldhgFtxRoMofeJNvaDDXh/l+usV5XuZ0+hXJkGUmNyjGCflYU0lZ8Wi+dPp3w5LkKQUXc5fpRJ/s
hIFKYq2a2seWPFf8b4fXiKxZ9WWjwrv8+B57mtZfxhSG0EahfUzFxWYkJtdA/G5+JJjHQluRKULW
p+SECE+5dcc00hpdM/XG15Skg/1x5ZKZwPjGHOnp4PH2VAZttaIhYdk9+ts2wamqBEqXegaUduis
gnSSxOHdWCPXm0S2xYsCNIt4AFgY3otUoanfCjqrhAFFE72tz80F2ahIAmNCqJBoWSK+S4LgKNuu
asMb3CDvXhEcQWim5si6Q73ULdJnKa/hnaDFlc1viW9d7UogK2xFYj89xcuVwYesPPRUfPz9jPiC
ADEoAjzsaxOYO0IVj0lRnocDqu5f57ZKqJu1N9NiP4gIDKgHPd9e4R1pFsaYZNtaXqd1hu1W5usa
etmwh+gDAfe4RT4v4nB5bPxNlq6R+oKZteAZfWnn3ZqRPFqGZIeJu6m0+lQgvu4swtvhf5qxXslg
RLrXmlPBx1AtkylktttbI4xEk7jI8grnEF4N9ZTpIY4SXix5QKP8t8oQQI7WXg1a/zV3UnuX1FAy
g8Ec2rp4SKA22dRfLFy+rij/TURJxUhYel25UP7asf7b8yd9unJUvFyQQuH+ATejIrxBNb71mHAb
jNOqrjF46NleM9syk72vxFJtEs6rfdfUNqqa55FYOv1Qaqt4K62DXthO/P02KxSs4A30gZJgnbVZ
NvZ1rlXooPcZYFyP3WV+8hk1zZUGyF7Mt8Z2Be+FCiGPqQm2AuJohiBELq2ETfVYrlTNueevAPuK
ubzZbckmCaW3RVBTzMbXd6DUcOSEocaPKU6J5+6sSqeR7HHYz0c12DnY6bmeGiFb0hC7x78JCDub
k90XksO/TMUoRNm1WWTzXnAw9ZMrA2IT/i9CNtqtki5n9PRNlpM/eN3Oiu/NJaYJYxhIli6QPuzO
6s6faEaen5yXUVnQV7xcYjJ2nTfVV0ouVnkfh9f9rd3ZQyzvuEN5ylK3BrQYUxC3nIIwBoCKw3q3
B4iiEf8ggu//vBuphm10EqO3kjneL+IOhIYjYh5lHDz0qL001QPME9aE0Nh6jvPxGQSd+UlupUV8
VEnPXjKbCTJj6UZ3Ltau5WDjpsrtR3atGt6ldCjRWaLeEvfqMmkuTn1Y85NTp1fa8oiMcfSOlLdY
uTZ7e+Zowb58bp5FFAP+jxrusXZoz73VADNgZrWY8W/yApxh2BwPfKYZZljbRstrPfcRu0u3owEO
oylcnmQE/ak1oGz3RyHpsLLmHwSNh0hF9Wqe9OG39wpvpn3aPCE1SkDv6M/FPe/Qi9rNuNRYVPlj
10AVdHgt9cx6STRgK4gyikoFSVB3I5sBDxFoWdYURscfynGWx1p1pJaUURceU55iVuTZVlFMvZb9
JooEMxvqKhS4x2TqGLe2uC5JB7ffDrNRDIEvmQwnkXYBuvmZwVrU5s0gI/SYlI+w5Dz4Fkw/cajB
TogB4ibWLW8m/8DpYF+26/1HcCNlrqhFWukJYtwZAPKufXPfUSxbVkrW42Y4sgQxttR7yAMye4Gh
KA83aBKrDB0UaFzH/I773iJP4xH5WbOUfxJL+VD0e9LtrkZ2tpmqGlLnkMyHOgNuI7I3RW45cOeh
Y+vKeRgrSDZIJZ2KhIV64UfniNRlNTk28A4tYfFGPDIsJBDKQoo78d2SKVtX6qvX/5R0FFgLK03a
w9B7jd7jvXiLzOF6H8QBF6RBZ/oWIvYiCNjLHTeqFH/8FUTU9PkmQFUMflftbiDUMcq7JE0zo9oo
NTIj5s4w5kK05DxjBPLHZaK4VwYfdOe3nv27ewR2SpEIO8iJNuJ816y0Qz5bSrD/oiu1Cv7BHv6Z
FYemf7pCDSD6ZTIujMj+W0qjJMVRVUfEWWoeh67UH6R8ofo1hCsMmMh6zP4qkjU=
`protect end_protected
