// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:37:12 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Zbi/UnJFMcOizT7g0hUgxeIlAiVryPT3pWz3OnxQE3c2A0l7XdAGucRrNMC+9QWo
7EFM4q5cmE71bv5U77HRmCsG0lpyo9EWjsb9AYihYaSMYQ/dJK+usBmLLkt1ELPX
5JA3/W/xsZiMg7aPOUJdm8R1FH5KuoME5D4aZ7r7Heo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11216)
H6HeYO4U8yG95UAXus4HYnTLTOaHAjWEWCyrjFlsddFNFJ66QikHxES4vYCBJ5Oy
58HwO4Tepn6IaHm70LjpQk3vjHteVW9nL+fL138a0Y+QDdiXyBTmLgjJcxigVoZQ
oI8yPdNOqVah/djEgKZsHVPyhmI8Gsqy3BaqKdXKcVkeSy34BRIcwiFNM8nJ6ybg
6dY+LtGDSq4L7s3ncypw6rBzMnNJwNB+uMHrG656NrejcJxKP5xaXo45SWXnNmtL
VObohx9eoNllIVmS/44fIcqGdfT1eQQ5O9GVBaWObVE7WlhdVzkrxxzNV1mHVAVg
NTbpdhi0nydbWFFalKs7KD/obA6ZFOQBHHjRUDaXNfpT/Z6Ka2ohGkRa9J/TKjaL
VTmHkfN01uDeyR5xElSDlz1KCmo7b6PLUtJRuOxY3tzLcXn3SeLwZYRqVGaRrm3f
B7HlxneQj9xB+MItDNoUknZFiK9JhPii1jfFfCACGJS7qHc4bvRpFyMNP+1wvb7B
7zXAHwnC/c/AYtIqKuMnR2K5BaneuGFH23BrHNVSqwRwGkz5mscQrD0ScVFgCsrf
DqUP419UQTrjFFwEyARoZo4hjFkWngaVnhSQy3pgW/G+3RUjl0Krfcm8gGTSWIFt
rTRpG/LbYsTlYhcA5qh8K/NpGs594GkaNL+Ob7J+Sx1HUFu2KFNbXrNjBQmDRSlD
TFysf7u2cV1KTl6PfU2xeo+nz63pfq+866kTqvAz7Q4UyCXBhnlqaB/KiWhi9+0P
IeO/JY/b1ErSt0A2Tukntfl0qgXxnqJjuOYIBJ9nAlYvjMCoF+hZvb9fNFs6aFNm
vl2/eJyWGvtLeSykocHsQViVwHLJV8jfkznySfhZOAoMqbzGchUpxuy+KJGef9xY
cHE4OOa3CXANYHnvMXeSYQ9oyMZzNEMRmR88sgKmUXCRF35GWaaboJH1VPAHDiZz
9WGmEZ0/L7wjkhq5FCypiSEGp7opb5R26d7fNlH0EpKAK0Xo/EPUr2D0Y1bIWcGD
/IA2fyUsBaMTf7pyGKoxzZnX1kQIn0bw0TdXiO9YBZnRYqSaw4l4WtnWEkqU4J3u
5KQBmIiZ347yc0Kj92RHTPaxGWzbxR8oUZnPGKiIb1Fi/gJ8Bsz6Z2EQ4C7QQ9Xk
mbTc0PK6WEzWcm6YD1IRrrexIUkso/ZJJmSg5/eO5PHPV5ZvnPLjvLBQwoxt8umK
i/w4YS7LzX52gQih78P5FVWyLGdtsAAIwKTqN+5ZNMDVkTAk2eVeS1vuIcNOJq9F
zxg6xSQH3lKL2PSZdqvC5zRBwHDjFOAsYo8NY/peZNnBRxlv9gS2WxvY3UNFZ8Wx
rs0HyeenLMwDlUz/CetQdeiFlYnjN1b73zPCYcmsGfL637Bd8lWAEEmJUQ+leB98
5ko/K0CWjbv7+zeJP7xanPQnoysaVsauLIHDMrG1V2/01+nnolWJSxvpbQS7YMqf
ZWc6rI1YXXZ6/JUoCKJdx/0NFz+/bZ/DkGB+I9N45mQd076PQYTMKgvlremg62aN
jpeNiasBRuRbkbfBFReCx9J8AL+B6+gQuMEHbcbrdGJTKOiap3Po7Wh+9+QPu2sF
IzCset9sGH1fJiwjE23Y65QyN23ciwAjz4dvWElp+wULyUJGyzMKIl63zoBVQOF1
Nh76OhRk02YBYOQ1GGZnQ1F0LCe+dTA3EyVWj1/91i3oRaia0LwacKYlyAT5Qo8K
YZU+W7IDtJH1ZcP7ziJUV4BoAE7Qq8Y+cpM4VlTKgfJ6vX3Ad8aU/dGuaPFRGQ2W
IlnCc3yBbIhlie9Dg9B1cZMHFIBhnaVafJinY5/Ovb8geA/EkZUTcs+K9vbZ9rDS
KObnD9WAnUBNoBNZC3Y9gc3a/5uHyKuD2b3RSmp0ZJ+Soti3+95vDsOSd9CQuwMF
T+IycLcFM7066ssRiPDu7WL2ceqLoYGTFgcfI15s3HL2HhVsuM8YNS+UPf4vIxh8
lrdaFty74tN/na9awNhq5AJJfP/1aldN0iOOu1aqXXOuDKq0ixM+wlOtcptJuym4
7Aj3VAtLpjKxFLyPhH9+J2j7o0h9yuvNMRA+Mqdb116C+qKHv0Ulm9kG1cYouNJL
r3RIxJbEg4HniSSq2Xk9wJQmb2TFBSfHJb8Yh+eWTcDE3OYBbNJlK9ODun92dvoP
OIslbYbLVwFOuf/2lejML1Hk5CxHAaKB6QGnkqVeVufh31OrtWJYzQQ+IPvxV37a
OthwQmK9ZaBgUTEzgQKA8qjmllf/j66DCxKiArKHD7Cm4GN5qecYYm67KLEokAWI
Xk5Kdt1qdZ6ar2E6n5pmCNPTU97MX6QYRV1wzItHXE5dLpKMdNlUJ1us5Jrw7ouq
wc1m2GRqA6JRifCnCMRaZa/uI0c/BOalyEbB+YCMX0sU3etInJZbyfiia54ozhbX
3j/n79Q6HG1C1w9U6LRprRXGfsefDzdkR84ucA4YqvEt9+S7+wVaT13hAeVqc6j2
RjVmzL/Co+n43QK9farzpFqCBZ+NfgqTPdOgMGGZfaWyXLhTAH3EZHd+tCDcuKYL
ntMMPlyG9S7zhT6/kQR9Ug066Ke0rmAx/PUw2uK9nLR6aIXKhT2hEq9XXFXhfK8h
I3AxpHIMFq1WxmrQq6Xy5sOg3GjFeT17NmO+UCCNkdZ+zRhbDRVqw+7ZXWVD82vk
kghuyhvKlMGewFpLzC7s5D0r1VBkwGjFIe8R6f5UilDEMHQF160P1VOF8Ax3/Mr+
QgqVLE3HeNN+T+RhIUyF3OM9xGjzpV6ilOAmJwEl5sDBUn1ECaS2yajBS96WqCE4
U9uVZzDxLJXO9/sBtugbI7u6IY1Z0SOn5wmInUg6knkZXVglfsYLOjeghm9ijRPl
9tjwSP7YfY7FxiJ0k0m7MA/QxrXOsHZLIg5Db/eraYfGlRHlZP76yeGalWAKph74
/yD8Pd98nrAD4w0Y6j8/PeSFgFyCFZCt4BM1P4Uzk6/vG278WGt+TAit1RYdRlZR
jpZA2z31wAbIKQGBrl2LeayVDoLoKnzP5H9JGzixMQjStzEojLfLQJHTgxqTl4dv
/DMUtZARq0bElVGKmTf6YMebA5/qxaKmnyySmphPbBcL8Rhmpq1S3njjQ/DEzYUY
ApqNg9JEBdPcVa3uPtKJcUP2z7DEwRl4nLOyUA6vkWO7t2G7gPrjQQdu5mZEt2AB
e0cHHJCsvC9Wf12an7zgoAq2G7Y97WfUkiQttkmZfI1LhAAdb0NvAox0HP1Zmoi2
PI4EfEtC005f4bfQqwbJZVdTYSd2EVoYaDhrBVGTGU698Hulu6xb9SZxyHdHNXyD
MixaaFxlwEmoIsCH8T18FrhjV/kUMxxOhb7Romh5Q4ZFJ4rkcM7/bAKrPGPB+sNv
zCOYUolcY6Hd0nqAxSi6Kkbhe1ONxH+qkuVrp5JS+gnVsuWEFrGOsOWaRpHZPv9Z
sKYhcrikE1I1tKLrkYAlKFrjX9Vfn3SNpk67K2IGkGtvIDIq3cAVFmMXEbo/qAeg
qTzl4BzRcs5gw9Ebsa9vNvjtB7SRYkZ5ss3rL0mHYVzrBkbW71NtpCu//LmsYFEf
DkSWYEB8N5F474CdgJY0C0oggfQpAnZ/mzraRI5H+KyCEnMd64IE76orKEyuAKeJ
fgA9AxcgxQC/ueWWZE254/qOUbIyKJdmNB4qtBpBvQ8etHTnTpq2QhIXgGh09vu8
rolo4t/QnsrNsY+HNudWA94YZNODiNDElV53wsPc4dGo81NpgmqkYjFuVajlx/j5
rYpSAbEvB2YQLDEWveYWCRscl0TfT/KFfzvfa2rAqqBPZ7bcvfpPXvLKduhrP8e4
G5n/9m/+PQCcld9bxhYKJ7JRkWvkPB2OqPhHXT5/DD34MBSloDCCIpyrLYk25aEm
IRWVcu0J4QgBUXiNvukgw3PueOA4Te2OMlhTmIKLhCiJrczV5Z98JdWRuMh9uzt8
CYcL34JqurJU0k31+SkTX/4kdvVZa57ZG4mmpOrFeBRa+Rk/YYX5NoZo1btBoGWT
uo09TyGTL3Z+uBG8E0BUS2x9uAfDdTY0NeBQjJVoJ48RMpWpaQ7xwRZ27Ombjpwd
5Gmm2VWeb3Y28YLdPEBTrWptctVtYTcnn2B+68mCiwegnwLOywjkoMxfqfYwGQO2
HRxigG+e6oIsi6KlKpdpfIY+OVHB64LSq+Bq7yjuVPxkfhogYQpa+r+XJBM9f3II
Pc0TcqfWwJaShk2+FqPUnsak/IBD1axytV1i5OxiXAQ8YxiIOJioDMHGaSDzNKvp
gqoPk1wdAnDKdCEe0uy6wwoEHt55p3DAI/tfTzRcU16R8u0toUyzNUd7Yl9aMiYq
fu0OKoIN5KHVDGmtI4pNzgN1QKK/WEZQw6l9MPobTBHP8iZUZcp2NWlF0CizasAw
lNRjlGTfh3zWq22eaTqhpYY/3H6RR70vcCCLol02CItNxuLlQhzCOHS8f+7PMt2z
GsW6A6x9S43nCg34HxlSyKLKe42H6EStw5yNUUw6we2zTLgSPTg93SFeaW64fnF/
GtDNfxZquooCebORph09W0hWqPOEX501WXBvY9FC4GysvHl+9SFVSnnnPWqK9zWc
DOTy3Gkm3nonahR1Ofq5Zd5nnICGVttEY32JlZcP43M+axKLs8TCda8tdtGJfwMo
xsXdT+fwqBChzTY4A79zcN65vlAGsv9OKjTgS4zOTckhdsiCQ2DyLzzRJk+0bbu6
QmRzm1BJ9F6N3WdT2y1mCQkwxExoVNCW9L+u2NlfxkBFhdvBL9D4GrVTgFoVCsfo
bPt//qDpQUzgAUC5c5PAG5veVgbP0cWrXTZQQ/WoG4mU6IpEHLocZuKH+Hszu73i
jwg6MSN5Sc3DLo5sFR0IQAuZO3k75u0XGYCEA3HVAjdqxwh3/lzlIC7UBVPlopXc
XqraYXb0IT+MjBry0l9c2bIwPC38FRHY1HntsrZEVyeS40OP2su9RhOjea3UXawX
aWqL5pvexu02/k/nWHkuuk/dyanxI8xS/vqQNMLU60mYZG6PsCvZs92UlIJSrFhs
HVeI3FbZkpftxN/BHuf/zuoTILrPou2gggQPemyViJCJeCmXx9AWIrUrW/7gPTvg
FG9OSxtQjDaB9uVrF4xfd0ot7t2O7GKjdi2+NF2Ok+wJk1mF91/WfHcjGmJvN974
JV8zZHZsei8m7ZlTVqbULIDBCWLVD8JEUadXoV0N/4gJ1nxwWMnRDIv2RcMqya3n
ZYoCqlOFnkj347/gAH2x3mlmKXBhJ2ztgbVJG8v3cloT5xjVESxPD9+MGaXfqulB
yKAZmnSvRxNdIGyN4ehq1LxcaVEMlD3P+ysOkKuQvB/55ZwCzbP+nKHvs4G9i/Vn
I0K5pf2fVRJi4zKomneH0qmWhyvBVm8JB5ytFo26uktW/kJFaTsMM1HbR+wYVGxa
tm7m+WfJXCmCKEdGSwZO98ZZERdhqbD0rlNQlU4z0ceKYwvkbqriSLMwodGDRbfp
LDtL3JrCOc1MawObQ+DEt1A+pTbqMExZNUkOfHSObXeSL1jpEs4UPX0+fxIxWKcI
6o7WaGhVErlmrXj1F+6W5K78jApl7vvYavDIJ4E2lZyQJgROCjE1piYKv5K4JI8+
aCWCiJwvIYcfu7aF79rh8QAJcvRUSc2LGnPuqMHg4aDAERWMsYk1o39s/+Xb/oOY
pRBFwmI4Mdn3VoIO+gSZCZ07nC3cz6XzTGvPGSVDrxb1S+voALsvAZFtltRaniK8
i2WfIc75hceYzcz5lv6csD0C/C03memPGLGu5MHxtiKG2w6rnUaoHfThBmjd1JnN
F/IFJX2tfIo0VPa5S1cC8SFNkcuu9WNe4nPDpHMfuE4GECSHHD7/kLayqJ8RRMBb
GJ1/MzLFuneLKcVnoEWjCHLnnmtf6pWKrO5mjD9QqXTlsoi/CPyEuVpujf/qQLHT
CXV1ztRc2tjO1jrVdsCnDu3v9wZPELX4mbrjP+UF8pWZL/s88HOfcVRv7La2txN3
zAy5mPUEvdTwDjgnEfTzapA5HgJGIeaSjOmAPu/5bTZ42rqrKu0CevCdnAz84aOc
KY7R4T6hePwkNMAJ6hH/EfoHV2JNVgK1GBWNIl6KqHF+hRqAkQcusjOc4IHrMkgY
su4JeKDr2DvS3W0TkJy3bK9fcZJxUhCYA/IPYrca8VPSosFMUbdCoKBnSWx2h+Wb
JKJIFavSpxAsWxZ8I2p/IerAohpZnyfctXh+XcjKPLPLIRN3qdoklbR0QbRUlX0c
UMND/2ubmWVi79pm0fj88SvR48koKkryaGaZQGFEycdrHGyNqtYVl71GHEIDBmOE
dkligDyt76zgAf/MAdjw4ETjcw0Prv54A9NddW0YglFJmsAvwnoN2JcJiDC9OdhC
zKVkdk7deYndDqezaM5aIzkE9O+RQ/EAS7HE63suKE0ABPbBOmVHrBhXbDReidWo
evBBplHMlmHCaAYbXLVhwOt8kWOhi8aSBfmWgqzu9ZOBBnIPBLUDLnSduejsc4h7
/jjJiS4WdRcBFiVE3TEyHAbqy4FYxyDI8TkV4na9MgJuDYHpEgE0LAEpwDIbqvF+
jmZ05EXFKoE7zIJM8OWBTLddpsPop9aZX9qazgPvOjqmS8V8R9OcfFXaCM8lcrJU
SCq50NiChL06gqNQzqCGhGpTCZ1LTk7BW6z8UfQyiJm04WcGn2DbOBfOnz9zfkps
sck5hJ3si+3u4KiEGGWyyYxoQ8i3NWzMQoKD70v7M+glGKSyfpBCkV9x6gG+8hwc
41nJeKh4u6mjN0ZM+tjQFGC/0ln6Q9s/8cMWtpyFhGMQ4ZQfT/pXU64ixpKZX79U
Em7lWQHlOkl7x8m46snt/3iX/ZhkGIVfdGgQLjLHRToG3Lum6WyUOkuXgw1sbjD9
7PsyXlWzOFHmYhoD40EGlCB2Ex5KeLo+Jr5mKKmTiI2zvIA4SldamUKKuTCbot8B
eDQx/BQ1Ur4cFiGI4mLNsWTd/fO7Aa4R5L9YSN7Jae6YI/oaxcgFGc/zEgozAro7
FzpNanNMPgk0v1v4qayo6fNfsFt42M8MnPz96KVxp9vPhr34/6r/5ijJPeiIprJB
IWfDyPodx3IfFvWeGCB+XqXI7hWmwE4noUfV0IuEop/uKfZ2SAhY7c8QITF1PU3o
KHsJmtMh8hXL61IJEvROk/PX860lkz8iqj8C30/LILmxv4K2pnCaQczsudgzZYhW
hkwWun92Ecn09jNcYgvbdQqO4ROs2S6T/UW60OrBsv4NDJ5DbQKHy7H0Sl1LVEpQ
dqRzMququN2qAL4cinkAug0gJWliqYTMrO3iqLKG9Z89pbPfD2o2g1pJ7AV201bZ
XP0q8qZZ76SDO3B59Rg4gKnvmPgowB6JrLKdKUVgzV8wBQCaOsBRkAIx4d4olhDf
IsdbSsWVZG0zMuYwCwqRT8f26MXYt3aEqatmITcQbK50miOWusPn1OGCvwJ2SySK
mYXaXSLakcYPs53szr+EKJHC9dLkbNuzSpjKMR+jZpnYLnijsDU6rhw4X17YVOak
nMv2xphzEzru8nhSuxbPZP1QHym2yqaL9I4wASv+UlWX3vhqHpaPU8G1zUhi8yY9
jq5vEGmzkC8dX8Jh3d6dUNEca5rFmrIH7slNgwuI0L/BW3xCcTCXEPBAi3StZ4DZ
5b7xVQC9lrCwVlL4evTkyv0VqxjzK3uEXwvkXQV1Lv6K0XVwtlBfoGAHvzKyqreP
CVtNfbiG6NIjfadm8v+BJEGDkNaM+eKX8aZB51yNo9FJS+OHaiw0+SDZKAbf5Y4z
rmz9lF8f3PsjmGqiOtSS3MMHJhBxf3k+kDKVCeq/nWo22ETjmZtTUueb5q8SeZo/
SD4nhCV+Oa1WgB81P+LBu9hIcYAysts06di6S+aEN9yrDwl+LRO+J5bfApFjO2FZ
iRa6lTjccjKnSMNMnAGyPpSv5GXbwahE6WnepLnyw8oESUj7V920epfmw8IwpK2c
m1cunzabM48SmnTt4fzHNPA+4YJUGwaxu96t/HA6aMFFy2KDnBR//06umMarqfFM
nm6xd9U1Q4nW2f7P9UjsYvvpeDk9aHda8MjBeiwr7JF5z+X6E93S4YPP2GEh43mR
9J7z+Jy9PZx0CrZW/kwkLqS0dPyUThRaNxVFsB5GYSBlse66RBpmRmLAvxoDMma2
6W2oloznlxEc1ooEPhgRB4CyTuQXojZsTWKDjEu6QK2ySwmK8jDTqZouvQv5Egd1
36ZKh7RiALVuybvenjdcm1keMcZ9Fpo14AYeSoDlORhzq1vb/4QcCMEJArwp8aAM
34oK2bP61xpr/nmaPHaUtq0eN1JxZZ+IyAMEG3BDO3QvW/oKiym8wgmGtevXDPtm
Uv6C06ji5smpGd7gAOpK5lHY5jhLlIL9G7lpLnAkF7kfCy71VjeMTBLOj7f+4WXF
C2KT4q8n6srjlRM7rBrg7eR4R8ZRz4cMINh0UJOkWa00LHr+3Zn0UiVXAWA6Y7VD
v5fpA6imPhE0FaBDW8/pxuFjZ+pW3AXdE3jju/S9yjYf2gBP1rdi8TOMHPWZyoH5
Cn+sI63t9MJpsURAE10JrKEzsN6q/OlnIRFm7OiNWMKetf2JRET+/VOdjiSZeqn+
BsOILA6ljQkw+qM9U6mlO0lkJ1G+RlI6YBHvQCNpUgCjo53ZCdxnJ0FuMqlP81ke
wIHyo1en66DQ0uo3EHwGaL09z4yTUGFevSc5S5fOVzKcs60yUjUMr/mezEGFcr07
3dMlayyKJPfIjDLsZCwX+OfrI5z9lBz+qRsYtjdlGnxkPD+ywINT1jQBfCuHh1RM
EGa7a7Jjdvp9AWTXkxR6lGGI+uaLiQZF+aXD8vpEaeHO5Y/2Hmgu+Y3FbwtL8wgX
7lEtnIR7LA4iJ3osHyjUSe6E+NOt/U6d4//lfGUNWbiBklhxrthJ6VNpoHsXatdZ
XObB9cpGcr3i4IW0ADnn0lYdGQIMCiNTbtjmcugMMkZZoB8p5d0K/p5SuHWocdV0
lHI20eN17FvptSjdDxMHuIYJfMqgN5Ucdvf8tNzpL8Xzjt8o/UEM3SU1b5sQK03W
iROQgE4GoBQyHxQpKps/PF5iy9t2JSZ8jA6dWB2DPjIYnjq4O2kWGAnPhEWlqJR7
9P21UPG6t+DzSYNsFFDvwLgWHuN4kD4NNOzGubjlkyqSMyvWm8ksDeMaDg0AoQGu
pD3Ofqn+KdzRBTrl3RQLyfJEgwZg9WNj4UbWb8d0yh5CgKmooqg1PLPWwOrItgu4
K3jVCOmLYfM8NGWVzTEelz5xtzLto8PW4X1/Zur9jiZeLOJstil6wYpZ6s9OmcIs
ElFNWhsc8eDKKpBZ3fzI5pAerqf9noylg1dLlu/bUf2gKARHnXi1H6Tg5wOTwzj+
6+c9E74t3tNUJz+3U35LsY+Fgbem2xZEy86c+PKb2vK9O11TfH7Ha2vpHA79BMVi
dvaMJaPlxgzQEYHZYew07qmZFlDEIpPsrAazGNF8wveGBwXgs1/pKEcbkzUqS5yZ
M5C8B+4UwRFpolKTJjVB6E/va8n1/ejK2rwUL070PzWvg6IfnORyAjFugNCs4Oa5
mdygf8pLd1RrlDpEFtGe2+69WztRXKcMCAZtfNid8x5zcsHu3e6hnx8H/hiEfY9e
189tn3fdgRL8R/Dfj5zSKUP/yI1F8GgZSi8xn4q5Q+ZlnZ5/xm4uP5VARz9a46E9
uXMQVRqr2zHAYTSB9B1ZvKUD7KkGwkhrX49rrZLhs0wJEw9WWYhIlG8w0NMX0a5N
rJX7XstvlLEvSYPwtjLYyRg+dysrB4sZCKZV0uiFNeo1AtM3uiHuQ/C2wyIW+FTA
a4i/EYOrnm4zpJ7gdzxUxoms64STZoB/NXRAGcYu/ZfUNJqqgDtIPOXxEKQoKKAz
CZ1O6w94YkTpN0RVhgsz0CeTwJ/iThsAvs2JzE6LIn5LvEryCPclkr2yUCKHuQoV
2t2tBEWMv7f0rBjhecPni4+hBhAKUd1GJoT0JXd1M1n+gbVAndK8xvM2Cb7xnNCD
81TQn4po6zLz0OSMHGeUvNL29E8Ro0LBS7Kbbco6h/Eyzev1x1IIws34znfNlvPs
UyYQmDmRVzi4HoeeJbdp/LjCa0jw8PvhmeX5nnbIXfMZA3gtdaJGtd50EN/vLMAr
gX2cgQQrpMHpSxfH0HqBnWDO23v9qY9LMlumQ2TXpsiDj8laK82T1Jeu3FCdi9oQ
6Z3ZWbE4FPZZFmuBPf48ast2apdi1bwRzIvK3pk5qTx9EPmDCYyYm6aSZyPPyLqF
yhxCi7QI9Pyd9eAStLHeH5CbI/uwikN+yJx7DZ7+Ci+BbER1+PROslBMlpNP4Cn9
HASAVSqL8CVyn3hniU4KHIYPEdWzPzxugyjPEHdaS0z3x2PE6ZecbVRDZ6DDeyrD
KkkRPWstX55jImypp5NoiMDXdTtQTTUzvy0rhUbwIi6GhvQIZ0wgxOUEUDtrCroT
ZUxVcjjIbQNXLGo3KmXfZxDasZ/Icg9EkvGXy9aTr49p0OGVcwATP5fBQ5LIm7i3
W1jp9RV191Pbbw54850vZvVQRubJYGUN6BO5ynVMX/XIK3RE2GoM2PRSOZ9ALbeb
lsZlh9S1mX+uJs9/btWuRDBc1+eNwm9/Tww+zpfZYhmxqZk9jl7xsSDrlFRwdFUc
nhP82nPQM37qNFJPwRBWVGa8RFehFFvCNvNuXvFT9BwICPJJWGFz70J50N7FwnEz
Ma1fAq4c9pONJXoEtw1LzlmnOAVcUKkIyX5Yo7t9cs4z/CDRgFjyEaDjRw9n2t5f
P7L6P01iBufaPNBfDK4OvsoCqBcRSc83JvR/UJ0NjuRnfASKOdzwkjSbukHbDuF0
myqvSDqe1dwzqB6u16j8p5ON8L37yW/GeQEPt5QzDP6x7hVETw69AT9FDNX5wnmd
QGGnMLeJ/c02VAk95hX7DyDcvT0hbkLnxd77zwaNU13uOsPZ31cLTeWuRkX9ebo7
NTpSka6ioJl9pcR4V1jfHRVLlQaBtGf0L7KVIax61LSxl0fbebObeizWHRQ6uLnA
OSlMdUzQDVY+kyqIbCWa0cnl2uN3So4yCngw3N0lgr6K5bEgEliROVwlL9u2j0hf
VyAzZonKxnTcKHuphJsfQz7mRx8sS1WQLFlHseZY3YbgNsgkmri1hjgMz2jCvrvB
YdZP4UutYoA2oLG0kRAISdsE5sExYJsBGsD56lEy+aoOBvjxbYxcv8QhuaWbbztN
9nv/ZEbrtzx8RhSKUf+IVOrBUo9649Iuj6XsXQxViKL+F1i5F6ogkjbAR5QcRzVu
alrVTsNTrwgXai7NnbhRvuggz4pK8KNXNMO7XEIvnIHVNUZ/xuIUfmIfHZbJ28ln
mAllkjFH8FJVgt/Y/pxDbqnKQHaUaZZ/2xotvEbGYNCUSnSjmRvjOi6TiXvuCKtb
JV3/EYkxOAEoPTQctDQYJwQoY8BXPeyi9+KSq7ddwe2zu3uml2NeUs+k7AkAJ2Kj
b7KNN/Pic1kv6pRwYlBiaa6plmZ8e+84M654BctexzB2Cn33Gw2OuLv2mhS86+5L
uo5K0AGacSPoFCXuipa+oE82dUUQ7BQSl4ZlNmH2/MlIEOnlj04F97MFmadKiCEp
dPdSTyQuMZTS6kdR8CSHJNnwfU/M5Hgv16jpoXEVUdge0fFGw6oJmBM4NvUdnf1U
ksf2zEvP/Bpfpb2FAgVrR2x+7XS8SnquBis9GJncGJUhb/lnuMTxNT1Q70QS8XM4
Zl8vxKC9myyHD/JtsfkqzZPkD9DSSzUoaZ0nPfVRJaAQP9QXcXBlOKipmp/TTGH2
+1I2UsdMowgQLtua5Ckwsjb50mzzS34dvJkVDavrBZsuzeLsjQKiM1z81OCibSHA
hQhyGFPEx8Gc7EiVy6+cncfJaIPDAUb7fw2QL2cGOAUsyWpK3d6bNugvwglSIxyR
x0zMax7mIqtK9fnDTfnAZcjBjcECGwGGMSzLEKMWW33OskemnAoV0Eief/0z9J+p
JILzQRePoi9YX/dwMqHTR7oML8L7VupiBWCw/qI7Fa74aJKgQYdn8nXUess58Nps
gp70lazBf/qOxaXPJ3AsICpT+6jcu9JdcnxtzWJq5bHaihwbYJrquML9lmhBywIV
YkmSDqSvBKZllEpC0p8LKGUKJahnUjymq+Y7e/6ZPEbedg3/+Q7CHLCNitWyPZDh
vYe9m+Eu72fcW67uXzteKFFjmGLuNr3nYRDEMVQPqTISTFyBcoFW4J8r6TR4z52A
FIYuYTmoWJfAHoGP6uSDKA141sFSE2hp/HKiIq1eKJX+ELex7ThJfyOdrqUQs+2a
zWtjGTsVw77CQlcnrst+cXehRKyD9sClXnv2U1faiQ3ve7iji3QWurCqryigW0lq
zvhhCYuBDBXvF9cnsLemRxNJSYK8ZiiJF5MoJq9nSVIydX+U2VUKf44fVN2puoEG
DU5Qv44xqwJSlhjTPEOdSM6AZ3KtLrnb5y7oJQd/wXftvklpS2+OSWnhrNGXFi2D
rahWXz8ccf/N4hI61gdX2iGhTNs59ATcm637Jp6lSHxn3ZulPN8PRmlgYKFO2gC2
hrsEYpRsVeF3EuGB/FhisfOIfBcRjn08qLjQJRm5wWt869PDu+v4mldZgzaqSfIM
AsJHO3Cxzoe1Vok1wr78T79/S8yZGNsIM7YIax5o1Wjarx0tvI0knL6JBFZuh//C
aV5D0alYJJ2cOTm0kwFDSOGbYqAJnfOBRcaTY8/dSTChcHUNTpb1IzO2XM9v18lU
c1JnpAd6yPm1/d1SmG4etHH70zQSbFe/oS9baeY8JRtv9LCdWZ2FAF7k56N4+c7w
Ga7n91dI6BIrUwItApIZFfErZsEG8fCHSoro3qoMx8H6zEnQ4LtszNGQx+8anrhl
T6KoEOIcx+EXBTG9oP4dXLfdoyQxTsX3BYOlL+djENtDUiT/EZJilyDVOew3hq8d
rDNcJNwMXUFiVAxfW9ewZTceuNbqISFzDv5vBRNFvEppcZpUwrBfCTzOwj+T+OA0
AnHhSNLrt89xIgC28bpeGEWYRgVwPY2ky8I6bo0AEDMgL3o2dWewcKFALxoDakhQ
0mkCkbKvs3VFSBUvJOpuzoW0Y8SrWFpFGEIQLE0rz4agsaUuIeoHhy2l2yK6I7AN
43JsJ+oC8Q1RoJ1FIIdshtwD8giGSpi8pJOVBYTAnTolSh2JtudRxEmGZv0HWy6B
LEKNnKUgevFVCJX2MpE+0Xj7ZdEvQ0TrIDdgnZ5dRlIKtP+yCw0hzz8wjzCd8cV0
tH0rRu5C6vmwfs5IK4aRswHojfcJf68I1/1m4yb0WZ18sDbsO+lhS+K8JbNUUf5B
ozjqhyFf9MlFaRjTOSFNlEDh62YDjZyCsFG+3skUuH9VoXVcvyXRvX0MP56aYIfN
CkoisPx/BviPWMiO4uGGmyNsQ4xXN7zmtJayZ+Ty7YOyFq4mmpHvunspyn5J0VWI
h67ly4Frq2/X22V1Y2pWyqNbAnGbqsdjeuALhwiVV4XTdsQTqd53Iq822J1kpkuQ
wpWqErnyaeu/IDwqom+5hiquINTH9cEMSrZjbvaUkJ7jWK2FLMm2g6ED2snH9DuP
2fVG48b96ra1uXmqKjGVfMI99exCfKueji4oLhHL+pVR0V4FXzBxYN4S7j25E+ep
+CJypO0+x4dzEAXGLwABXJcr/7tWrb1Tl+w2XqkRFPZtm1k3TH9BC+JU0Uvfuxfl
PsGNFRr+HdN6Xo+kj8NbhMT16bnJZ0EZOIaaH5S6wSaKRIMuIyX9dAHRfB8Su1aN
pDOb7zIEgrwIgW3XpClMK3D2nAxvMQaRs7A5iugeVT8ujxBN6/SyACZ8aHGLqajY
ls2JotOt13H+DoDubOQV2JQqF9nEpExRKfYy/rfRcjYzC8GFlrN8tOhQ83CNlL5j
Nz2lI3JGjd7oL3T+t9icUYy9A7UPLpWp10Timgb2mAVcF3nMQoBVtzrbId4+CH8D
XLFaAaE5XWughsX46/NvwxKCcHpyyUibp7GGBZ+h+c0TLti8A5GKYxsgKWfwaqWX
2l1Y1uv77YNx6RXeod97keSh7tJVW3vlLTbMggYbPzQfOHZ+bhsa6xqUYELj1nc+
CjMPIG6nhlueVdHzpgddjqZjIYTCAwaIiZSmNF/YrdShgKDzXfA6CJqLP7eQmBXX
GihcnSePp6yBsf0HTkJnV5F0Uq02HqiKmqezcz6ZzCZutKXu8KLd3XzHOwJekvDL
02710zZT8x1jo024waCFllFPoUT/Eewbllqjtf3Nl9Bp0mHNCncnscPWag9GXJDu
/9iFz81ls5nHBN9wrc0D2Vd3k9f5sDvSqDjP46CF4ARV3x8o0BJphKezn1/WhdVu
3Rte5yGRnsoa/c92DTz9pixVyUNKmGJ8ZETUB2U3FzQAItlY3bgRT6TZNdACsMJm
nsdzaRYfJsW40dWkZzu7cW5c5oac0pNWmV5jWtehu9tYLXSJBCFbYb+D8fnk8dpA
Y+e8WoZ48N9D3bo3vy8kkOc3jbp8P0pjXohJXsMAUwtmMSzg5PvSmOiAkGPXURHH
K1P1NqUiWS97aGPeEMzGH6bj//3NgKGyglFXCK3I1bHgdbNZRQWUPZRgyecEJQQY
Doh/Xya9HohYVFZu4IrR2vavvaLMtmGPxAnQI3xJ+0DbgT2gmU9SmyTDy4lNMuaf
Hwr0zn6tuS87wBhpT+8i/3VGCZfNrAzeoiJqyjT0h+8wfImDyvV2k2K5KQLu0KXL
2vy764knwsrLxtHSG6/xWxt1WhF57HMhh7HgWYp480RN8+3S1G7OHJwZsrKCPxKz
Tf481WX06DdJuGAfNbZKKZrWbQ/C/y2UML16qOtmeEHzmGrfxOADQaxH5Ibir1fa
ud03y4WLMKpPrDjGMaCkNPmZQyLo6bfMJCifMTvfftw=
`pragma protect end_protected
