-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
R7+Dim7ynROjpN9RAQRz/u8G+kjo+K3Xj19aAUfzqeLealCiiJpn7p1LL4VwThAoRlONUUQ3+0w5
4NiqjxnKbfN8Yk6ch0gjV5qUe2rbslOhpJY28epv3/HPRdyhGPDH5zOYi1kpCWSUrn24pOn3VIOh
Np6f/QzghZG08CkTXewHmwAAKTyVtgke0hwr2L8tIVFcMPsNU59RwfdqSJpq1662sK9cazBKKd4F
Kk3/qyhWjzSkH5YBQm44379b5tcmc5pJqZ5Pzwd8nFZEmHj63OpY6GNsXLtpsBTCcNVXocRKiyUU
Cwo5MLAr+ZikTqEwZITzAFl2izWuKzKUL1uWRg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1072)
`protect data_block
oSY/EzbLteTiIsUfEyMMoziwEPu2RAj2Ri8W1meG1sLGLaoMQh8ivbXGkHmXJf/q6wMC6Wy07lSk
exxgQgG3nCxchnQ4AGcixvzAXvrC+ZYrZ38odHpXAAJ7/luX58jHc8BNumsm5axUjRfityaLPTEB
ZWAhZ2bYSBDnr4EEb8lYb1LHFHTV1lO4/DQpI2gRNpF95M5KxgbWWfhkH3JcxQWbMW8EF9Rchacl
2DuRzEAEf4nCSASVQgKEX4iliFd+SHPZckeoBlVLUO1KUgzKb4IpCtkKH0tAprw2+fCATXIyTORW
tYgzg58T34/zSN5j00vam+OB9KUdwh+DjDVQQcJCvhNv8oyjbBBKO9iBTRqEJmaqFdR9uxxvypjo
Wf0r95YGu1kFt68m2WEj90yF1je9e5ZQ9tLLpFYO1PM3/3a9UfJP+RCLDSntGzRi8btFipRBV6Gp
higQ+3F2TpAmzst8ifjp8KjvtrJZI1xplzQCpEptGdLYW8ZyfioDjipinwxTgecfMtwtq5Fo9ums
vLAWCCJ2fKYxFzc8kYXIc+8lICQcdjjnpwcry3hxdNcXcW52+W2LiJlTtmBTzGpy5Z6tg0abt8dp
5dqqG8+ljrcM8teQp8kRk114vrRPAlnLiBezfag0zJhNSXsuqjsYNkxo2ic8jQ5MkdIg4rybrp5l
As7JnUmA1fCy1kYyvRbQEQ7VEvYRRfmqK5C0KRZpUXYgTandPzh1AALilYCzA6j6yJ3PPm4p4sNc
jyqs6O5zjJsfs4aCtCv5mtVGZk7i2s8puEp3n5tpbRuBxPvQn6mvfPVhcbnYgxVqTZSjEn30AIIm
Bsx1+PtaBuWX7OJ3XCtvNALuOB3BTaDemkrRwaadsM3SVVMC9P9uO25rK2iOk3K8ffO00LlCRfUI
3Ca5giS5Y7zs2tcxqSLvI5A0eYqLIb8dNP+O/E70SneL1/juL969+e2kP93hyCnasqlLZzAdQLhN
ADGTFl8dEOwPizWOa3j/xRDysR38GMXwaTucQWTYN+dIMlCHoF/n8Zivr3R0iQ6ChBrzyfODjI9k
9jP/aLargkdRIEpODXiT1y7FQwLP9QOp7e9OzD36bi2xWgGfAcCXb7tz96PxuEbyG7pPvv+T+vAL
o31j4AYm9hyjPPEZpFp1krCN/FN6W6dFxKy+YxD0QXJGBgm77Gdyxx2hnPn5XfAj22xusJUFrIuQ
xM2HP4JyX3aBnPWF0NHfP4iCEYX+sZBQ6trumVZoD14/DyLymzsrEuRo91T46ZCSjhkxH2Y8z/AZ
FUHAM4wNnAypnVLUe9TYWX4TG1IL2j/hn3kr+3KfiVa4rJ9M/DCBxXgIDCLBkrh4hmosqVnRdyYS
hdW9K53WVM16Hcg8I9YWedOfCiqaLnOiHfKZuM8aNCMkZOcuvKY04BkmsRW6hw==
`protect end_protected
