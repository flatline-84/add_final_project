-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
czBhtukrvKqwoc8dElt1X6OS1g4HjcNHpsg0dJjL3+MUCzbTwy7Ud5sBmq9Eb8NbEuNnSAhkvPt4
6BdFDItM+FRVM7ISS6qHnbRoIAoVdL6vsFilMpXAwp6MuNsHdr0A6QPGjhJfUgBta5JH57qWRY7K
Dpyf1p9H9patbiBVxUImwi0WQQtI7ri/oL7jl39G1JS2/vxsFDACK2Tq5b4cbQSTY3Z3s3hpfcgb
FM42AFck1HtnxztHpqBeKcxbv9p1KAjPyt0Y283rlH7/yW5uWOioWhvTEN8mfqKm7QNSujHo+TCE
o86F8C3/3g4QTIKAPhAM6rRpmbzlLm2B2NVaug==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11888)
`protect data_block
dKlq7i9Hldi97/5xDv5Ul6VRFBDycxPpz9XDS1GdRGRDX0wqJznsb+GnhnBlVY9HAED7gDwkeyf5
+VUTndnIOvVrgc5Fxv3/15XfgO0XekrkatkWeusoxVyObWeHd3kWRR8aUt8rYm8DJsXZ5Rh/oKpv
emT9F7TteMZ6fNCFdAa7CYV8a8TEuPEZw6S1bXyTALbsrmaaTokdEX5RfL7rDXqXCnaLKPrsLKaZ
90UAS8WuJYBIyKB/WCr/PPtM55MupHbKt1auQ+WJ03NmXz1ng8O9Je+nq8NJVh0iKefiYK899tJK
xv6Nca6xBu3Z3rS3oyO0h80xKa8fDlpzU4Y3nNMuUCFbk8jKWrJBfc+ALVSXuDsUlDiVeFwdX2pA
mOvgccFNo+f0klTZTaMCRF/zTuNf86BRLyuPNOHw7s5AMv0Z6YPGe/qtk+mTIiH6apqQmITg9Qou
cC30L4GKvpyGeUzCzvifnpe/f2WHf2PBGvLJwZIkYF5hKYMkzw85mgFLYNRfR5cRrItaIUQ265LJ
C5bWkVSqQQovZpGoDR0A8eLIM/x+9dWG6Y14q2DvQN+a43aWdDfMRDHG/QtXDiOi0pTjoCI3RRnF
JBWt8ew5X4gjPIzIxK6ebTRmeoseY4ZzvdnHbDelM9RT94d23XDs/tbQpyqSl3LwedtUQBWz7Ban
dz3rgRfhT6wRp+0AAcmh9gbDFy+pihdeUNnnFEDuJDPYQbG3AGM/X3zIxB6Q50XBNyOJynOsUdKk
0IAkDHEInEFWBb5K0Ptn5Y7t0ZUHZA0FbzPYzTYKGiYGYv9t0SpQKjHPnT0WcZbd65XnKJ5r+7og
UJCcvNw38CRNiejcCy6Z9TJEL1ToTBuBSnl7Etf5umRyKTvk/ALHa8xn71u4Q03/0H21tXTI6ryA
na2k6YFopNS8kOO17Mmf910MGnMl3YMvzLqPD9yW9Ueqzi0Y/7OeS+kwQOY6RUIZfFks3iQ7FbWP
hIX8eGIzsChJGRJ0lx97A0RmAPpuThxw45FNzej6OciXNVJ9poEbEME9LYlUFgeaOCCd8yFsZFbH
OL13FS88+ZES8kJ6xDGMEyNBRFLJ4Hegg2xf3Mw2W/UGB4LZkLp/OkeY70HxW8+H11pBY8R6wX4J
CR/jMz5ovtNgXMaxEhNQ5PQSul5tJMrdCeM7HmGQFlQPqk2i5V+hdlciNw5KkxbCBz+4rYI2AO0b
6FjfYQjCi5wV/gzCmCiculqS3zE9021ds84nbHd0n31KQF0HTRE/3XBGptHpzCc7HPw7GdO2jmQh
xv6NB+HXEiTRd9SMm+8l50wXX0VwYlxZQjPli/9a+hoShZtiOZCZ34JqaSJ9d3zuC+FzznpbNEj2
3brl1+8ikn/8dfKyMlfHuCGWSEI9f+ChuQirdlIMaHOv6Rix7xbDRsZ06LHQNKFb3F5WrLqh4UVF
cMdBTM/BZapVZzj3fwaCbTk2t/B+fh4H5MOQaEMJ9Whl5fIS8PZRSpC/bjztqgANXjzT+HI5M6kK
K2TEgXgabBii6lZcBjgvM2E4eMpMGKtE5WtsRluTDa7rdavtZcrT1tGJrv3lAuRh8AXU8yvMT/Fx
h15GP68MCRC3+G5urYwFkkMjRSqDbIYRs/GJ12hIR6MAcVufwwWdrLPDWMWidXlZmSY3NIcLZlEK
Sv0Yg8BpbHFVsbVMrXyVL5pNlj2rXcK+shIzdxT2122TOvQix4qGzxAy6SXSEcsGNAQkyRqOlEoq
NDM4loe5KJEpJ3irTScUTB5vDUiObx5yH/Gm/Y070by0kISkuR1HcTX5CzgYpz+0rAahWuP/+iV5
JIGHLxlYMXpNxHhpk9AwFDhSoWNysX3Y25HIzrqV4K1fStVbLAzydC9FNVRf0YbjKnOPXjNml/gC
NpEIws79TBfcy3Aa6WZ52YECqAwskaBlEoz4Tr/+cyfZAvyjskwOkpoQwIAweuuVmFuO1kRbqZ57
dOVvv7J0f2g7MDm3uI9V5a3QomMyjjC3DxJnUq/boyq8mT6Lz7nxZpVGrqveP72+enZnIpZAoWUC
3tKc/DCIzwBaKSCF8EbTFDTxlQl7hPTL4F+1Mv3XLCUFcdCVSOqxP0y5WP7V3plAGJOArKoEwCMl
GsEm6rm/6Cxh083LmTicPizdSCO0u8WUwlCdYknwYgCByV0ZwgnCCLh2HcqAyrzubxkrOVmd9wy7
F1mnPXNrmciv2UNlGmZXYJvrR83gS5CjlG2LMqW0NAzhSFU+oMYQDqkczgFHjtAzq7PtyuNyp1Zs
EXc+Mw94g8lFS5OBYtxhvb+5XaAIG7iI6V1VCQl7pVM/f8Q4Pu3lwBFA6Lu+mi2XGwhi3wcoIUOI
4JaDjLNrzXosAD4cQmhXiVdaUHk8HJQ4faV1hSp0mpD8YDD9JcDBydYabDP/ckwkFZa7ik+Aghn6
X9/kfTSZmE/XjyedmCu0sMwsJiOGMjiFIN8GkLDZzYVW3+MEfLX92wtLrQUGL7Mla52gCxOGynjT
+epJ8IooQaLZlmIzzWRxjlHMF3G2MrTnusgH7LEekWsGuYGHi7yGHCvtZXWt/TEFJTxZnlqfq+/W
h9EViuTR/QL/tLmDF2F56XYm9DkttCp4gIvJ88X6kaNa1E0iDGT4tHhv4RcpFV8Vz+4SHoU59DGV
K1r8mFRl4mM6x08Pi1SUWzqaTwjgl2ajosnHWtXrXQKNx/fq9pRLGPKz7cwiywcl5TeZ8H0T9G3C
LS/HDFo1/B5QE3RZU9sPmH5XTFC8gBRgS38Uc5jPSTZlU6AA2XGtWY4Vy9Z4vqiHSe9VbhgYXZ3x
FY9B8rvyOlP7QJBra+9BVvUozErgYUipPwRZXMnRkMw2fN2pTki3T1DbRCvj7ss0vkASx1rjCA5P
xY3VnoHbgNif+V1aw1iI7IUybzb4LGkooJkRLwipaxLpqB0mQ/rNx3mdFrraCTLFzmrlbS0t86fE
b9YvhhR9LG7X64FlpEeZN3JBFpGxsM+AL0CtFrMtYFy7Eyk+pP4Bwe6aqWS0Srj+crCgKt0n34fX
FO8RU5nDjUBHAxk2gs7LDPL8FUV8/mL3TUmBgNl/mMSVsqgQA4XQncmrG1hOgtK0coc3VTiCg0Se
3EFn+Lvac84w3M4VaJuCl9XzSn2alR6LXyKSxyA9a9Y/H9RGMG6Pj6gKAAGBf+a0ilBj5HljLRyo
1GuQ3h1Ws/tP/PXwmWMOjb4J6n2UimV9kIOnwJgppJqat/26hn4OUHBy0c6ntoWIkiIY7TQKBDZc
PF+K+0RtvFnBVcJZEa1hE5ztviertMg9U4sodYPjtNzYTK1/NaULk6yYL/6+CM9AYTJ4qX53AYxD
M73ytZnckCJLHMSuYvA6x/y6WF4xqVv9N7/cGqnbFmUMsT3v7Pq6jO2qeGtu/6hLkzqDHdB2U3CV
pgBG7eSMhsz8uy0QlF6yZyPKHBopQVHWSoBhGNlkutPHMGx0VVPvzwwp74w0pkCGkAggvVee4hyl
Ivl29wF+0LU/IXZ4CcMjtXtcdkzx8lwhRBemAgYDBGl1Y2ID47ee9OoxGO2gvyx9WFZQy1WOwqHR
u4cJd5PKTSPGcuVsEpikh+YaAscdBAmieKtY+Ws45n5zcFOduDhTIc8Kqv2Kjc0OCN+ETOSnlONN
1Ql8Uwuym1uAs8XbCNywrYpdF3NjX0eHTzQCy8RWXl8O3IQ9M8cfz4TWncJEe0YhSg+aG92S6A0+
S84zB7AXaIoLBCFuvOJ4UXx8IGJPPJrfvCFdA378So8i8lWhk9wc/n5k9GS+6DFhyAebgC5QbXrQ
QqFKoVmUhVjMElt0XfGCEDqWs053oycMlQs2uNpb0bbsBDZ4n+EquQHPLz6ThzRb83+2yMQCMWNo
KDe7LeKB7h09CNe1+RNWXJV/Z2TfO+Qt7t0TBEALfhS9xST4iEyFI+vs5RDbiL+6JdapNt2nReEp
MnCo33z/4DlAAMkkIOmyb1dpysl6BJsagzrFzwFD39+NWSTR48n7YykfNJ6lsqZK9VUIdosxPslq
BiceJUYSGKFQDKN42o3792cAZrKEsVHHObsjLUwNwQtRvWx6Vjda2dMQqwvfUI42TZsbcyQzeThU
wdp4z0bgRIs9O545k0qElHA4S/sjBv641CwpNVrbwUlpBTlOlnDP+bJL3XZckV2ag8LhtROS4Te7
+zFnBNKjOPaW8Qau7WM5oC+rMg93JRaDCk0K4fUv3syGa2YUIfNWeO2nsEAlb6Wk98xDw6T7/YKk
l4YCiImPuWcMSHctmtYcTCgpKbl1PXmegWGLL72rMOotT6rKWtfXsB84cOM07z6XBtXjcSHkZkOC
fL/iaoidKHNnxC3q4m9VPqy3wPaiX9f2BizvS6+sBzCdX/alAtWM2nAAYi+4fqO/LxEMeFUpXGZr
J1yTrWp7Azl/Ji6Qy0tqeidHznqNP7eMviJ4HFIL3mJSlqvSJeNXj0q8MZhTaq3Jkzq+sshgBsrC
iONGneQUvUf6MQJNnWJLIfS5y8pSU9ty0dy3je0+jf9tLLCbkhMy3C2VsqGsov8mYHM9d4j+YNey
wTuRTZxni4wPW5juk8vsvnTqXgSUOaMaDcELEI4JvB93oQSjO55lTPtNXFMlKgQrLDq5jILROvdC
qPJWOf/EcrWKeOK+TpFp9hM88VZv0xdJ+n3ctPmwXLcGcrhZyRg+FjjVoRceDm65ZV6YgqZmgmWr
fDPdbjsi03ETGEoccZt0+mW+YkDVA4bxa8XFvEgPBmG0uJKz/EeQKULVXEwt8+vGj3mKP8YTHv+h
VToDE15rnMsjkqEl2I58XPKhct8cRV/FCdLWWKkmQprSsHs2LADZKqp6RES6syzcc76+BtNvmi1w
WLQny4kXbkxDMR15341PN7u/EDy/VbzM0EyOVjDY0hcAyv7oB0baaOe53k8hBKhv44xgURbJqC3U
KlEEQVFFPQsrnns3g3RJnXBVyOGuEo4m63sNPiA9gBjIwVV9Z7WHblHzf0fd94TgDo2npaMfk6aU
i+5hkuOgxsoG1+noK6Hywm5U3pzaUMj6E2iJH3b2vKrxbR647m8/TPt0pUqWK1SmkuoKsbj6En14
fG1FrgbAP1+KWHNh2rdxn5mYEO7OkeoS1SLpM03WcrZTgCIeEETlgSq0MlhWfzILnq3EYZ0T+f3x
RzpcxNLHtqS+yw3CHrJ3S6VNZqfO/MRpr3riGXy0gxChlKtYpw0uAm9lCx94ekQppw+EcXvsKg4R
ycv4k+0jmnp07j53AZ5P+IUsp+ywGnJk5D1Qu1vDymgkAbhPGyaAdA/lhtrSkPM2Ff1yUmy3Qj0k
DYlN+Dq4Tok2hP8HlbGZSJSOL6tspNwjzvu4QUYxu0+pJ4masH0AmqJArMi0KEumyIDw//DfqB8o
I3NUqqNGNF+lVpshYfxUnWn5w5oq/KWK6RJHz5d0EFddYYkLkojhsQcGjQpd+Sev0SNPGrTuyMG2
pwMCdog+wUwnVUfqwS9zNPlYz/Am6tvxA0jV8oGZLXvYAyMSiDldilyMQNQ9h+lrEgoi0g59DKMn
Bf++UhOqnEgabWbz1LwlBtQd6a4ykwEENPMIw4usBbQ4Aj6mU4o4qUrnvzVkuVyeRjPI/1d0Lpsm
YFdtbwfJOlb1earEugt1/sA2NzylG6/IAumiotInkcFSeo13R8XDBDyAYw9AhLLNy1c5lAGXoH19
ADj+jHG/GzKJZV+8SMj2+aZW+fVwr+Uf2qRX6mvZuQc3qdB+7eD12Rrh2NkMkVQEGPdsk9bQim+m
wZx2hpkywzqdirRIHhVCwzYNQT0qgZjPxbPGslo9OxPjL8HM24TcDVE4OqCJwr5NDOWvnQTbhNxk
KeQ0cKwVk/Mc1oIe7c0sT4AvB6ZBz9/GQa0jXL5DOimvo2coHxGqXV+jbxiqI4XuFNU9q1f+89Sa
8L6pnAgFjC1ksoQIXf0yErhR1Yr5cWR+zFEyczvu23CyL2eNP+dUMBoOzObfLwI3X2ZuzhJs6VXs
seE18rVLwZ9FZokDmk6PsAfB8otUrXTPt5WnvcJhF+AZLAk1SDw0MTU3uxr++yp50vFgWsrntmz5
RpLk+ksLSSf3C04przFENkCw2qCBOypsz7COTf83ALAm2+rHCuicztnlTmiGfZaUJzmRIKufPpjB
78gABXE4WY2BrYmaPhscLezqTIeADErrm8w1xm/YLqBKBhz+SGqxndB47x0jPwyY8nM7unmD4WtC
hAYb8/14ZH0CYpkDyJ6FFan78mHvT0RJ3iUAYKzsBmWXrDESXiCqoA59xV72Dzozt1+B85d2MHBc
P9ejhAumQPA+erSNUZ5ut3Za3Fuk+EHjAfP8tWFKrqIuMdpejRJaFeXIzcDVIghRjJVasMtpHFtD
t+sdw+eH/rxLxs5L388OpwqI6iojMN93XL0EAeJLh4kRDulvrYBXj9R7CFNYf5vizr4xVtI9xS5w
+Glmcv5RTRpFTcs/O+sZgmKYXDdLGwFNGTGCPmgs8B5uH9VtH6LVonQWuLfXoUUT+HVPbmSsMwev
F8Pf3elgnmemj0hp41lMDnDemok+mCZ1pb35eurZg6VpFYcg9IIMkXtP3IBmMfCxQ3+SNwJDbJDq
H8FLWkMScuk5yNsgoVeC/TlFayriUcEZWTVd570GLa19Po9XuYLxD7OnXS66KdcZsIgGZtsl458a
pRY+OH9BRGUGI2A/G1WUzdAVXveXl9dNo8ykIdUzbiWXUVok1XV5PuI13nm5uzAN2NGtl/KcYk7D
zp0pKN0lknA28I9p0fzIyletm+v7fE1+caS0bodr7S16XwQk9DaIlK2myVyhuak3XRaJA+7QI1wD
Sh5drbwFmQpLAQ0bX6Bkb7T3206eaKNf1g37Rx/2qLKj/KDh1JSuv4PmiQzloCBZ3dHc2ioQ7qRZ
NwsJvFxfDlMxS/P2midJ1GdJ2VP+fbNK8GDm1UvtlxzDvlGaKFzdnCsw5N4peS2xhWu3fKIz0rg8
hvBfAWEe0TETVVslGaC3m5x3qd76tb1bYcjYsRE7maCRzLxvX2qe0VaExM0H7fnf5mWFZVHN9dHY
2Dq9Kq+IoqsuvP/CLl8xkb9873wJHUVTMUUwF+bAnv4A8Gqgol1Hob4rMi29sX/IJNCeXAVpuXJR
/E7ZFdrfEzrP48L5DlcWHn4MyEWxQymzZmjxYh+d8v57nTV0I2jtJLkbI1FXKK4U//xbGLuHC6wh
cyB1q7jqBKFXQSmZFC9aVSw1RZT9BbCso5DlEmWAUgvml2NwM/5S3Xfh38c3zTO5ZIN/fHHW++Wc
xwmnitSHsKDgCakAojSOmbppm5k8xbqXJHYeZjrFFmnsbPJz62EGXAzqw9xRSwZQvNVxum5sD2XB
iGo4wiQhSbjv/EAakSF+j2GiBpu1m1/z4jWPw+uog1dLGcUEtG//2gB0mP8SZmNfsKduX084eq1K
cn1ePumIkEeRQMybApdeAShYuzlxkkZQwjt6P8UDlDQfPDHZ0Tpo11DBHLOzsIp3ETUOOqiy4iZw
5c001bxsVBXPsidVwA5nUa0v8+2esb+5heZ5jd9yRndAC4GNnyKs8Ml//PqnpvfpPI7hVePKreGA
GgS7kP8gYiAgFalSfocpdaGVR4/hN0Bm7igp2ftZ3tlXvILWjSTswcgpOjYeQDsUy9saz4Gy08In
ty6cJY9GUKEgZkvRQXaYOdU334gg5KykfgQqjAytXSZ903lcY6ZafXnc3S93p8cM/OzTXgUWzbjo
XwwqsPe6+5Jdnfufamfdy3v2wHISOC/PO50/wBta4z9UPGxGnAe4fMiOce03Bswn4k0TUccRfx/v
YPvr5tH4ebSxIQ4nzIoqcmygcYXoxbMn9qmxhruZ+EYVJohjiWUMECCbarxY5i/WOWKPCh14j2jR
aQZHnrBe3ECoujmuyM3MUMq7QMPPE6ZPeb/cSPCA+LdDPYDakOhM8zOyR1aKLRvUO3+KWqAMPat/
XsOIdEQa8WfxQbmV85Z29cEvaSeLfsVkRtEzKvuy2rFR6zdTSIxTCUTyVsrqpy7cJWzIL8oqxk1Q
/txKGAkAC6QjCQRkdww0EUBz3/y5anV+YwVkmeE5B2u5P1//d5LR2tXqGrI0AZ4jlYT82fYUIYYj
o18s/NFQEigjiZgQDRtQgmDQJhheOjeB9bU94sKFbX/qP50c+KrYSIaB+jWKSn7MWiMcOgtvT2hj
QJH7GwhZrw6ypPli/acKA/sR+2DWBYNh3m/Y8FLeAMgln8L0NV7+ekoNCSZ9i1vHONsTsJ/EqUfW
BGtaVZnTyDnPjKzz2GD6NQ9Gvm7Jto1sSKnx5POHgvJkAVIkVWe7FmAQ2edjcyk4ITR9oDSy2wCi
iwkwoX1Td0zlBQ6oBUo7Am1x2IW60Z82Z0bC3oqkpyB9Xq5ua/sU1NXf25fsMMdMI+sqDNhH7rXC
XmHJgp2e2mjMCTTSCjinXvd6OVlDSHiAeMMEvEsjLfcb3pHhh3HJCwatg5A0TO1ZNhFf07PHifFu
kdeRP0Q5YC8YIVeYQoMpSFd0us5vqA4eR6sEpK7EUhlRW7vvcU3nuQ53twnQadW0ocpF25en6d8z
Cg3DfplrG73me4RSlZq5CtDCeE/x5GnJpTMtXsyUz5Q3t4ArVYPSFjyC7PvSHgQAnQ0PmGN90hbW
Hn+0voN6VmRbNIE2lVqz6JjOCsM6u1czhy5DEGpgvbIAWpSj4pZUFnHy/BNPtQzIAu7OwokMVGnb
piPOs+pNp714NHqnGkWbDWVx7MYpR3bokoFpYKkRRn1nszLkZBNGVJS0y2lc/QpKGqHWgxWDPCNg
W3OPr4iJudCdQ4YEiOWegoAE3PuAi6elcMM36Q43FR8SZ/fdcuQbaEzajvKFVRewR6qe28DboSGw
V3qOXTaA5N2gM7E8gqtfAHiwFqXlpi3CUgZKYmgvWju9WgnS0HYv6Ho3F+UbK8dPT/poBXenygJ0
hqfNnOvf5MbWpHW9RooDMhuy7xdERK5XQrJSRpQZVeEXJ9g3Ci4cAWvBLJ9Jk6gVIaO/VKEFgVyQ
s/qSdywzTA4pGjOa7I1FjQgfjSTm1GsMd/n6VdPxwMkCIsJt7HbpfL8mzTtJrO3Ls7KqLSOJmxdF
MsooFpLVWU8+/tv0N/iAnkmxzCRDX6ddfWPzkTSHWSmz5ONYjeIhmSl2hcSdy4epPCUiehDx9DF/
lwtR2bBD0aD6sFAmoktKuqtHs52uhuVDG7iCIy5rNEXW3WK3irEqOAph5ebRXdmkZHGY+17jeeqL
ey0NJdV/byv4eVpJ7E/YS460KC6VVFKVLkQ4wQhJOBjq/2tT/nG68hrV2dv3ypsDU+OPFa4EEHCS
oxWppzrR8N+O2sx4ERhu3aCPWOvndx1ez+sRurt+RSCvLcVCwEhA8jKUJVRhJaNsRr3cSmWCV70J
qh+UDkLAK6bCPySkIsHXbPGgL+k+YMgQ6Lycq+mQnfKCILX5JVeEvmseRRWoGuSkSpMUouw/6FFx
IglQJDPhrSSJ5kRkEb6s6a2t3QaCIhMoBKLLvpddM1mW5c3NZ1u4n0xxED34BcUCF3sUvUcpfcd7
wfJ2yQyfttcsUDOQqcE2zRqR5o7brGtxtHN26ZDgBbW5pSi9yt4yDgM0w/f+hAkzce6AQbd9LycH
2mRVm4cDXBcpMsa1q8WABagU5i0ujDBBF4fYj9YBeIK6cuhSGpbhCF9ujZEIfWyXHlw1HE1jWrn5
1iTZr2qG2uoSLR0ffeSG8ulEFz/DLnEpeNyEGuE4u17RblJx6/Kk6iO+T6RDjb5+14msuA56ccT+
NNAO3mU56ICyWVWU0hbXW62qHjXz1ulharZVFbFOvQhdhUOFmD1dtjwgn3LB/kQXE+JGLPRa5bqK
lOJpdaFGe8uO55Ln+MEnIy1j5oqSzVU7nFnfC5mjWJAcmTMH1UEW7mB5ymHE6HTGhQzT/Bf9MW3c
qhzu6JRRIjk+j8lpnx3c/77QiYDWnkFOCdqJQT1FN9tPN+xEPYXNc0LTWtuDfICLhpDgNWSAF8Vm
vaMpqTcZybnvi/iGIwB/cXojUsZtlPUdBxV8kr6BCv7udBUzP0alpvqyxV8iq65ygnBdxbU5gJqC
2sGGdrUyuZihMoKx9vdusaQW91zjYm+DJY+YAm0Yqk4vaO+rddeLPRNPR5E0+8h2jFDczpalHaRP
pyWStYVVqgmhcFbrBMxNUIC4Iw9XVuycmzi/V6YV09YpdeMEooOouWMH2xlXYJRbDA41AJqy9MQe
6n47dTlYihvkT6wkoM5o+7SktWwJxc49/EgCtE6mT8RQJgkuDmzeSG3ABo/vCcTTytcA6qI4lQGN
k+9f7ZuMwTBp83Sghup5nL2JiaP4vjGJblq4+ms12IVsspyBNdTgAOW8/p4O+Rie0EP0gb5Nj2Sb
EJ1fsqd0IcEaUURfU85N7/fyUaOe27lyONcjhzo7m61Gsw72kETCkceDm0d/tfhoemAc8PbvZrnF
95x9klzR3P6o4NZrZOt0XmrKml/RsodYMYzxhSu1/rlkkrE3BE82Gd+0CJECN6fgRnNfGja4sUZ8
K016aNtWzWXKyhjoLXGOptb6RBYOhO9g88dL9y+d2A8SKXl9jU2DfziwAVrQkwJy6rr+nL2bEU4I
RTPDVuA7+joWvgkKZGW2d6ZlZzdOFIZ6CaoTlUZmYUbS0pFpJTgQ4hoj8xa61O+FaqzFetJj6bLL
9ji2IYM66j5MfvXbcHupSRzyFGeGlgKHKV3mrayJtM4SK31LYMGV5s1Ex12m+qwKPbPiOnsjSiiK
zaR5ALatMJCmbbE7jpz9NJYN6IaYFx9RM8pjdO/kheaufWVUT2Df4eOrH6GWVZGotQjhNTx7joSX
N7v0QJ2XovgwJabwo2Bzh5uT16qLJ/SOWgypdiPaO+L7gTM7EkWdB4ei7V2qwPtmxDQUyrE+j0k6
4M+OWIhNKGinF1Tjn/MopUf21/Hu76PWAnrEDHyNbbPFQkD2PIe/trSjfllz3RD+zwJMO4/2QDIR
mhCPDZi6tHSQr/7cPKsCFY9FFgDeH0feN3aPSuSFUf4uNAsm2fQ6guDDh+A4ems9VhD3+K8WNRNS
BVwp11HtdAd/oRLVyGSkHPGahRD52NURzudSyCf7GPaDYXerC+DtyGtynusfK3G4AVUXAAFwVWt5
uV/waFW/P4Pgi4n5GBbCbXDtY9rc+/GiR2GvArjtKNWsb/YnlE14W45hyK+eqlJnrdAxgMkN2uem
VLNU/PDFNrIR+Vkfbkv73tlxzUjB8bm1qwrxYVyElzXvB5S2xmG6N0SpmHOXW9gAkbqRgQX4/AsG
+0mkfoJidD5YsQ/PBtlYwhvMDevz+JVdYtr5k3U7ODK5XWtC/3J3CQK+Mk5cPmlLHbzOxGfQ3nF9
6xpiyLQRgvCoaL1q0rYF5yqy5l1AJsxzNRiKdq9ejug8hAEBUCRVmJIDt13t6Y/4y959CjshqUOh
qFocI1kfCb3A1ROzNToRSvLhFDd9hn2gtgBTZRFQd4l4gQSM/52JvFi661lbtr5U5Bwy+hGJJ3ep
48YJn9pwA/cW7UsQ2yurMZzsbgbltuyvSnLJoTameF3zrE/CdWr/2Uc76pLdEJ/aglFgOHNIKkFG
iIHwJRXpOUzKJKPmYH7JQkEhiLn6Adc4oGlQII4sRExBOwrY9FsFT93g/Cg/95M19c2wgNX2DS0A
zawxP3E3UIqCwPblbqXzPPvbN1rlTmlU2GsRkDv3sFV+ZRJyZg0g/Ww8B1pdpeMmp7hqPKkZxLHB
dXS778usSZ87p+y8BnFIiHnplugm0m12ddFviSHORwP6WFHxG6hvhI4B3st3CX3FGhX06mfGluXM
6SJ0MPwP8KmJ9ocnyWuuDiXkk/4CvxNqPPA4R1rEr0GkfkvdtLe6/oCuZagq8ycx7+ww0wJhOKUo
nQVPUE1c+la22WsgtTUO4QAqjsLADSKPEk+OIt/yEuO2vX0Y+5wYkghZp7m+uDxwI2pNaibLW8cM
hcE/4Cr2IOQak6FBZs+1ShVfDwczYO0JX/61qkOh7qKC7cXdMUaVgBHfqVd9AVe4UKJAVsZHpiii
rEljHYjxPuSGaIwRr6t6yDuywAK1kBKxAhk09qo+PdA1D9bmzVYFEAOtyLbuUujyDg4WwuaRiG+G
urABubtOvq2Qv5JVKg3XdZhA7+hTSAtdDbTwm58n1y9YU4n0FH+lRtDMIV0VPQQp4j6jBR3WsxdM
qU4ounfzuS6t5kA95FXk6kbm33R4DxMpWYHalzMdFn/P6S2lcNL3W2gKEumPW0Z3lNERJ4Hmcb3a
tWQfzTQZV3lip2HtBPGGInB8NGPrkY3HkZCMYaHjgqeCr6hQwvVteMrL0o7blwOEbS9NkB5+bjhL
vacqjusqtxc+AIdOYYgESLTq/Z5OZrquSplf5uEnaza59wszS7mhc7ip4x3DLM0z9oCRmiJKT6kf
kW0HI0nvofbEgIHcUwoYbdRTB+VDMCyITEoannXtYvpdHEubW8IcY0Uzz8rvkNDUPpkOXGNxM1eZ
A6Dzdze4IvOprtZBJDTHsm/vvOOW4iwUw94zllObstv2VF4frCM5Llqvhua4odZtfJp3lsX8iSJJ
w3wd3p318f000SyDLf9DOwkv2nRBuFCB+BHQkNC/xu9aNvZs8OLb22n8AgQptHJoQx+LNWct74dS
QUIvQuLb+R289VIl9SvZ0FinoD526gKJhUwFx7GF+l9WuWt318xDkz/SUepXI9yg8Qniq9bto6bH
9xN0j1aqJWM4QqM33eGPvj9mtrpUeBxRChnT7syY1+v5ZvNtpnRMikG04nRJmbp7QuMBwntkUKjP
ML0lwYxYaRKe88Gfd+Vl6TGJ/FHi1gOefVnmMXScK2J03gUE2/ss1hVbQ0qphCFq1eK2Uo5V+kSz
wrIPZoZZYBQuvli4ch0z/JzdWY05+NopzrvHH/RLfzVbD5Ua/WvckphoaQmSwYPsWwm6HCf/51Ct
VXxRagwUNKtkxI7CzElSlw9Q6Wteom2N50MqSp39Jl2O9WG99YiYFUjhVHO50rGTRvWmwB0A09Ti
TsCZI8xZTgMDVJ+HOPua+WrDrfN1ZNu9JOc711ueug2poDgdxHVoShrs2dl6f8UX6k/kXQvLOREP
ZVjCFMLgh36Npw3D4BtGxfMWwu2p1QuriYUzdARgzcrZ0l3XDOxV0OBwM0b6cbWPY4LGVa9IVZc/
XQakZ9tu1lAVCIcCRAhrf7mOmnztx0ejkHoUx35pf+9s/d9GjQV0j435NMhqeTaPmPSNIRcS90f8
TD6De+UH2vJRkZQIJu9LgLKC6J9scapHgw3sezZbcHW/DwmyrUx/AFRBAxWlPoaJA1fSY+fV+mBO
odOYc2wJer3rsWDNFEozezWJOsizmdt8FZtusFrKZiiy3RmhaaXHDpF2vg+gsfv0kZRm95qbm0Lq
I8LwQp2vBxFw196M+iCi14BXwqAEzRv+5Tsi7QCuhISPqal3e6qMuW/HRxgaeWtTxFDsyPGb6LHp
RPgBiU8eP6GIWgfGv7FgchCOXzaAjYOEH7pohCqvS4RamYgJUN2vFLU+Yf2+QloH0tptQtJucosI
QTwym2K5yE7CR/w7OOvxuI6uiJrhYvT4AWmT3lFTgqNKXhXiij9UQ44ronQX0+yS0GYpq3XCG+JB
I0JYBdM7noLxHxn0etjYNvTaWjTRUBbfo05LEXXp9wrz6cr/WcwR8OJmTvLgpBvAoW6+0UMsy8Aa
Hz6edgpyJGXR7jOgSyzhDBgbPtlUK43Y6DZOJAAEib6cJv9LzeenBNQCBofMbZ1fZrJaLuUCm2Kh
Z89u0MIIT1qvqlRipM4BaUZWW2x5KwbKxIvV/QOc3i/dRJnQNqCCCoDQkyAWHs5k2HueV+FWTR8Y
t/xyyCzlit7yL7Br2Ax+CS0NnRL8xWM9At6RqQKS5KyttZ7ovSDZWYzdxBGoItVrEKRHcihP9PO7
8pSbR3qaR2CPk5fOxpukQjxCX0Jf3S+7CEt+fkcYIhCAY4CAxqlKOBSj+54q2jnR01EgDsY2nCKa
Qkk23+xeHTgzj2aAZr67srGFr0W81ON2RuvWuaYUSJS1qpcmY2k78kP9tiOxJyjXQphFJGPNXQQ0
VjqywQQJpNYuaecnrZyPrzYkVBh9xP4yojCPFQawdxnAuEeIUPuNpWzDMUYiTcq/klfKsryQ7L88
BLAXHm2HSVlOVZHkAWt5P20a8hvSnvsvmtOYd4e37ucap0f1Uz2ZdakADDu+oEe1LtimcTPQxSmR
56uVtNXZgJdUTO+YdEXKp7NwhUgl1tJ6OAkMxjlBQ94erUu1PCwwuCy3xV8WscbgJp5kE2mNwWhN
2brye/bQL8phi00mqI+s1x+8n8qaTRyXmtOOlCRA+02QNMgupPGgMhG4cfrP5nNovNQRhnkkijqn
NXEGM0V7eDIkOUcEQuNfBgNeoEZ67j+2KfHx+iea9W5aZM8O7kRU9OYgF3+kRyYkl1f8KRx4DLvL
kr7A7the7U11/esCIoEYmaQ2ssV7laFse4ILCzWRARZyS+Ak7yVDR0N/G80MVJ5GtVLjBj+hkj04
j/S269bGw5vRp7lnTXuoXOuQaHm7sfeIplDkldJ9WG2iZOD0edb6UiZHVSZ6owhFZP9BbCmWb423
OsmFtBguLAvka32/ocgHsSs1OCWpoQ/N56iYo983PJXgsAp8f34Evbiz7xsIPTIPc1VkWDMOC6lt
GEy8ASg2T/0crccw2A9I43hwH4wA4OHaIwrcUCSaON3JDM3ezajtFgx9L2YdQR72rwDtphCSCUuc
xXMeBhykhZsavLmqVNtao4+2zb5SsPYahtooj8RrgpI1ZO+AiMtBfstbGKvXXNX0H/dqnp/TCXAJ
T/9rt2EwVZ3df+Y95Gey9iKasKKxGg4EElbWqPicM+oOh3dB+qZWa/QZyo7ZW5xqrg8El4eluujR
KpayBEAzyRFcspKai0d7qu7DFKpwd7ZQRrAXCeu/l658qKw3SMMGMBzCwb1sVBYPKvGpTq0PGUnD
EkMtOb6U0Coc9V8v94UdOcY5dhFyD2U+vLMHYbUaxritiYV3ZSZV3lGR2SoC9Pn/tL/TJLDHmLQk
FH1tJdyy4Ecw5MNKJk2QFA785xdQ7G3IR30iXXIRXdUYZFs+rTBXUCM6KMbsnO6x+XeR1jeMEhmY
5+99cRwvRJ/1+metY1hGSh6wIFDwDWJxDgwE88PVxXEd0nBFWfa3kVXbCHkEYdavoCmg+zPQikf4
QJ2TCl4Ge5hpS3tNKoGVfjOLitA8BByKOzCSqUXojlbkx63nzFeqGTxofeuub4Bfo/Y1Q3xoqZol
VgyJDIXbH8k8vldWvz6icm+murNFOss6SW3QGjt8JwOwUQtpS2jQWh4wg8BavR9jvLyrhtFEeWqL
Ega6w7QH78XnMy6fPcsbfvFFj9DZAzWqsYff3hO2V8+GFnVSj9SVos5x2Lr9LzB48+DWzO5t6a5B
4a876sWvG2jvBzAYUfxPLxbhayANH/VHwVK6EQWLWBlZDeYrn+qQy/FcNaQiIDRMZFPtKH6JhFD+
wg7E4t6k+rFVGxxxqgYrsMtqYKcnpbsPIqa6piPhiF/A25GUXbjWXDX3Gb06kJ+JXQlRXDtsx5Qc
+L6HVsh+qBW22e/9nDrUpDNG1VB0mVp/P+lLeE/M17iuqr9N8EJz4UV+QNxsSYdOrmp/BIcmClHX
YHPp+b42qjI6F0cv76ttkCVa4ImK6fX7bxicROymLYqHP9i57YG1FEHsdvb8MM/dSjnX6ERJfjsR
uGU2SvLE2OQxsDA0orjgJBUar/Fnl6JwedaQyuu140M=
`protect end_protected
